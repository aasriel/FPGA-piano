// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Wed Aug 17 21:55:12 2022
//
// Verilog Description of module piano
//

module piano (sys_clk, rst_n, key, key_pa, key_state, pwm_out1, 
            pwm_out2) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(1[8:13])
    input sys_clk;   // d:/fpga_project/lattice_diamond/piano/piano.v(3[12:19])
    input rst_n;   // d:/fpga_project/lattice_diamond/piano/piano.v(4[9:14])
    input [14:0]key;   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    input key_pa;   // d:/fpga_project/lattice_diamond/piano/piano.v(6[9:15])
    input key_state;   // d:/fpga_project/lattice_diamond/piano/piano.v(7[9:18])
    output pwm_out1;   // d:/fpga_project/lattice_diamond/piano/piano.v(8[10:18])
    output pwm_out2;   // d:/fpga_project/lattice_diamond/piano/piano.v(9[10:18])
    
    wire sys_clk_c /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(3[12:19])
    wire clk /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    
    wire GND_net, VCC_net, rst_n_c, key_c_14, key_c_13, key_c_12, 
        key_c_11, key_c_10, key_c_9, key_c_8, key_c_7, key_c_6, 
        key_c_5, key_c_4, key_c_3, key_c_2, key_c_1, key_c_0, key_pa_c, 
        key_state_c, pwm_out1_c, pwm_out2_c;
    wire [14:0]key_value;   // d:/fpga_project/lattice_diamond/piano/piano.v(11[17:26])
    wire [14:0]key_flag;   // d:/fpga_project/lattice_diamond/piano/piano.v(12[17:25])
    
    wire key_state_value, key_state_flag, stat;
    wire [2:0]yinjie;   // d:/fpga_project/lattice_diamond/piano/piano.v(17[12:18])
    wire [31:0]cnt;   // d:/fpga_project/lattice_diamond/piano/piano.v(18[16:19])
    
    wire clk_beat;
    wire [4:0]beat;   // d:/fpga_project/lattice_diamond/piano/piano.v(20[12:16])
    wire [5:0]note;   // d:/fpga_project/lattice_diamond/piano/piano.v(21[12:16])
    wire [4:0]count_beat;   // d:/fpga_project/lattice_diamond/piano/piano.v(22[12:22])
    wire [7:0]count_note;   // d:/fpga_project/lattice_diamond/piano/piano.v(23[12:22])
    
    wire n73;
    wire [2:0]yinjie_2__N_1;
    
    wire n14, n17188, n92, n16773, clk_beat_N_126, n201;
    wire [5:0]note_5__N_45;
    wire [4:0]beat_4__N_40;
    
    wire n77;
    wire [4:0]rom2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(18[27:31])
    wire [11:0]data_out1;   // d:/fpga_project/lattice_diamond/piano/speaker.v(21[14:23])
    wire [11:0]data_out2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(22[17:26])
    
    wire n436, n444, n456, n464, n70, n3800, n3815, n3830;
    wire [4:0]rom1_4__N_338;
    
    wire n17218, n18774, n18773, n18772, n18771, n18770, n18845, 
        n5;
    wire [2:0]yinjie_box_2__N_394;
    
    wire n10972, n18769, n18768, en_1__N_194, n887, n891, n895, 
        n907, n911, n17250, n16909, n17235, n26, n25, n24, n23, 
        n22, n21, n20, n19, n18, n17, n16, n15, n14_adj_1435, 
        n17230, n17229, n17227;
    wire [12:0]PWM_in_12__N_452;
    
    wire n17226, n17225, n17224, n17223, n17222, n17136, n17221, 
        n17219, n17217, n17216, n17215, n17234, n17214, n17213, 
        n17212, n18763, n17211, n17209, n17207, n17206, n17204, 
        clk_N_168_enable_507, n58, n17203, n17202, n17201, n17200, 
        n17199, n17197, n17196, n15507, n18761, n18760, n18644, 
        n15506, clk_N_168_enable_512, n15505, n18758, n18606, n15504, 
        n18605, n17195, n17194, n15503, n15502, n26_adj_1436, n16860, 
        n17193, n17192, n16920, n17190, n15501, n37, n3759, n18757, 
        n18756, n34, n15500, n15499, n17189, n17187, n17186, n17184, 
        n17183, n17181, n17180, n18755, n18754, n17173, n17171, 
        n17170, n17169, n6, n17168, n17167, n17166, n17164, n17163, 
        n18616, n17158, n17157, n17155, n17154, n13027, n13024, 
        n17153, n22_adj_1437, n19_adj_1438, n17152, n17151, n17150, 
        n17148, n17147, n17145, n12259, n17144, n17143, n17142, 
        n17141, n15798, n15797, n15796, n15795, n15794, n15793, 
        n17140, n15792, n15791, n17138, n17137, n12156, n17135, 
        n15790, n15789, n15788, n15787, n15786, n15785, n15784, 
        n15783, n17132, n17131, n17130, n17129, n17128, n17127, 
        n16847, n17126, n16_adj_1439, n17124, n10337, n17123, n17121, 
        n17120, n17118, n17117, n17110, clk_N_168_enable_518, n13008, 
        n18615, n18614, n18613, n10403, n16959, n13;
    wire [17:0]CNT;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(12[15:18])
    wire [18:0]CNT_17__N_703;
    
    wire n7, n14_adj_1440, n18747, n10969, n17249, n247, n10968, 
        n262, n269, n312, n321, n331, n344, n351, n405, n406, 
        n407, n410, n414, n415, n417, n4689;
    wire [17:0]cycle_17__N_740;
    wire [17:0]cycle_17__N_663;
    
    wire n7_adj_1441, n9292, n22_adj_1442, n6_adj_1443, n22_adj_1444, 
        n5_adj_1445, n6_adj_1446, n46, n44, n5_adj_1447, n18842, 
        n7_adj_1448, n42, n41, n40, n8147, n38, n18737, n18736, 
        n15708, n18735, n9654, n8146, n30, n4, n18734, n26_adj_1449, 
        n25_adj_1450, n29, n16859, n15707, n15706, n15705, clk_N_168_enable_456, 
        n17139, n18730, n17208, n8, n17146, n18598, n6_adj_1451, 
        n18597, n18727, n18726, n18725, n18724, n4_adj_1452, n18722, 
        n18721, n18720, n18719, n18607;
    wire [15:0]fcw_r_15__N_495_adj_1720;
    
    wire n16888, n16876, n12983, n45, n44_adj_1453, n43, n42_adj_1454, 
        n41_adj_1455, n40_adj_1456, n39, n38_adj_1457, n18717, n16868, 
        n16865, n10160;
    wire [15:0]fcw_r_15__N_495_adj_1733;
    
    wire clk_N_168_enable_534, n18713, n10216, n16917, n17228, n18709, 
        n18708, n18707, n17205, n91, n18706, n17198, n17191, n29_adj_1458, 
        n22_adj_1459, n14_adj_1460, n18604, n11464, clk_N_168_enable_533, 
        n31, n9757, n18697, n18696, n18690, n10407, n10405, n17182, 
        n7_adj_1461, n18462, n18461, n38_adj_1462, n18460, n18459, 
        n18458, n18457, n22_adj_1463, n18685, n18612, n18444, n18443, 
        n18442, n18441, n17179, n18839, n18684, n18682, n22_adj_1464, 
        n29_adj_1465, n17165, n18680, n18679, n18850, n18847, n18846, 
        n14_adj_1466, n60, n18677, n18676, n18610, n17162, n37_adj_1467, 
        n38_adj_1468, n45_adj_1469, n18671, n18844, n53, n10074, 
        n18669, n18668, n18667, n18623, n19839, n7_adj_1470, n18843, 
        n18841, n17156, n18840, n18837, n14_adj_1471, n7_adj_1472, 
        n19846, n16854, n94, n3, n18308, n18307, n3_adj_1473, 
        n92_adj_1474, n78, n79, n80, n81, n82, n83, n84, n85, 
        n86, n87, n88, n89, n90, n91_adj_1475, n92_adj_1476, n93, 
        n94_adj_1477, n95, n98, n99, n100, n101, n102, n103, 
        n104, n105, n106, n107, n108, n109, n110, n111, n112, 
        n113, n114, n115, n18836, n8_adj_1478, n26_adj_1479, n27, 
        n28, n29_adj_1480, n30_adj_1481, n45_adj_1482, n18835, n38_adj_1483, 
        n16828, n22_adj_1484, n17005, n18655, n18620, n18619, n14_adj_1485, 
        n7_adj_1486, n8_adj_1487, n10, n6_adj_1488, n18654, n102_adj_1489, 
        n103_adj_1490, n104_adj_1491, n105_adj_1492, n106_adj_1493, 
        n107_adj_1494, n108_adj_1495, n109_adj_1496, n110_adj_1497, 
        n111_adj_1498, n112_adj_1499, n113_adj_1500, n114_adj_1501, 
        n115_adj_1502, n116, n117, n118, n119, n120, n121, n122, 
        n123, n124, n125, n126, n127, n128, n129, n130, n131, 
        n132, n133, n9, n17020, n7_adj_1503, n77_adj_1504, n70_adj_1505, 
        n17185, n9_adj_1506, n60_adj_1507, n18652, n53_adj_1508, n18651, 
        n18815, n18814, n109_adj_1509, n108_adj_1510, n18813, n18812, 
        n16869, n101_adj_1511, n18808, n18807, n17430, n18804, n18803, 
        n17149, n92_adj_1512, n16896, n18649, n18785, n18784, n18781, 
        n18779;
    
    VHI i2 (.Z(VCC_net));
    FD1S3AX clk_beat_75 (.D(clk_beat_N_126), .CK(clk_N_168), .Q(clk_beat));   // d:/fpga_project/lattice_diamond/piano/piano.v(232[7] 237[4])
    defparam clk_beat_75.GSR = "DISABLED";
    FD1P3AX note_i0 (.D(note_5__N_45[0]), .SP(clk_N_168_enable_456), .CK(clk_N_168), 
            .Q(note[0]));   // d:/fpga_project/lattice_diamond/piano/piano.v(255[7] 514[4])
    defparam note_i0.GSR = "DISABLED";
    CCU2D cnt_2220_add_4_23 (.A0(cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15793), .COUT(n15794), .S0(n112_adj_1499), .S1(n111_adj_1498));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_23.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_23.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_23.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_23.INJECT1_1 = "NO";
    CCU2D cnt_2220_add_4_21 (.A0(cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15792), .COUT(n15793), .S0(n114_adj_1501), .S1(n113_adj_1500));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_21.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_21.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_21.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_21.INJECT1_1 = "NO";
    FD1S3AY yinjie_i0 (.D(yinjie_2__N_1[0]), .CK(clk_N_168), .Q(yinjie[0])) /* synthesis lse_init_val=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(213[7] 218[5])
    defparam yinjie_i0.GSR = "ENABLED";
    FD1S3AX yinjie_i1 (.D(yinjie_2__N_1[1]), .CK(clk_N_168), .Q(yinjie[1])) /* synthesis lse_init_val=0 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(213[7] 218[5])
    defparam yinjie_i1.GSR = "ENABLED";
    FD1S3AX yinjie_i2 (.D(yinjie_2__N_1[2]), .CK(clk_N_168), .Q(yinjie[2])) /* synthesis lse_init_val=0 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(213[7] 218[5])
    defparam yinjie_i2.GSR = "ENABLED";
    CCU2D cnt_2220_add_4_19 (.A0(cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15791), .COUT(n15792), .S0(n116), .S1(n115_adj_1502));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_19.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_19.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_19.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_19.INJECT1_1 = "NO";
    CCU2D cnt_2220_add_4_17 (.A0(cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15790), .COUT(n15791), .S0(n118), .S1(n117));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_17.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_17.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_17.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_17.INJECT1_1 = "NO";
    FD1P3AX beat_i4 (.D(beat_4__N_40[4]), .SP(clk_N_168_enable_534), .CK(clk_N_168), 
            .Q(beat[4]));   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam beat_i4.GSR = "DISABLED";
    CCU2D cnt_2220_add_4_15 (.A0(cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15789), .COUT(n15790), .S0(n120), .S1(n119));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_15.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_15.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_15.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_15.INJECT1_1 = "NO";
    CCU2D cnt_2220_add_4_13 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15788), .COUT(n15789), .S0(n122), .S1(n121));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_13.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_13.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_13.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_13.INJECT1_1 = "NO";
    CCU2D cnt_2220_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15787), .COUT(n15788), .S0(n124), .S1(n123));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_11.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_11.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_11.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_11.INJECT1_1 = "NO";
    IB key_pad_10 (.I(key[10]), .O(key_c_10));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    CCU2D cnt_2220_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15786), 
          .COUT(n15787), .S0(n126), .S1(n125));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_9.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_9.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_9.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_9.INJECT1_1 = "NO";
    IB key_pad_9 (.I(key[9]), .O(key_c_9));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    speaker u_speaker (.GND_net(GND_net), .\PWM_in_12__N_452[2] (PWM_in_12__N_452[2]), 
            .\PWM_in_12__N_452[3] (PWM_in_12__N_452[3]), .\data_out1[0] (data_out1[0]), 
            .\data_out2[0] (data_out2[0]), .\PWM_in_12__N_452[1] (PWM_in_12__N_452[1]), 
            .n9292(n9292), .\rom1_4__N_338[0] (rom1_4__N_338[0]), .\rom2[0] (rom2[0]), 
            .clk_N_168(clk_N_168), .n19846(n19846), .\key_value[4] (key_value[4]), 
            .n28({n14_adj_1435, n15, n16, n17, n18, n19, n20, 
            n21, n22, n23, n24, n25, n26}), .stat(stat), .\yinjie_box_2__N_394[0] (yinjie_box_2__N_394[0]), 
            .\yinjie_box_2__N_394[1] (yinjie_box_2__N_394[1]), .\key_value[10] (key_value[10]), 
            .n18598(n18598), .n18597(n18597), .n18644(n18644), .\rom2[1] (rom2[1]), 
            .\rom2[3] (rom2[3]), .\key_value[5] (key_value[5]), .\key_value[1] (key_value[1]), 
            .\key_value[12] (key_value[12]), .\key_value[11] (key_value[11]), 
            .\key_flag[8] (key_flag[8]), .\key_flag[0] (key_flag[0]), .n5(n5_adj_1447), 
            .n18808(n18808), .\note[0] (note[0]), .\note[1] (note[1]), 
            .n18737(n18737), .n7(n7_adj_1470), .n18807(n18807), .n18803(n18803), 
            .n18307(n18307), .n6(n6_adj_1446), .n18610(n18610), .\cycle_17__N_663[17] (cycle_17__N_663[17]), 
            .n18719(n18719), .n911(n911), .n907(n907), .n895(n895), 
            .n18677(n18677), .n887(n887), .n891(n891), .n18713(n18713), 
            .n456(n456), .n444(n444), .n11464(n11464), .n18676(n18676), 
            .n436(n436), .n18679(n18679), .n5_adj_11(n5_adj_1445), .\key_flag[9] (key_flag[9]), 
            .\key_flag[10] (key_flag[10]), .\note[4] (note[4]), .\note[3] (note[3]), 
            .\note[2] (note[2]), .n18747(n18747), .n18754(n18754), .\key_flag[1] (key_flag[1]), 
            .\key_flag[2] (key_flag[2]), .n18722(n18722), .n12156(n12156), 
            .n18724(n18724), .n18720(n18720), .n18813(n18813), .n6_adj_12(n6_adj_1443), 
            .n18763(n18763), .n18761(n18761), .n16917(n16917), .n9654(n9654), 
            .n16909(n16909), .n10160(n10160), .n406(n406), .n18755(n18755), 
            .n18667(n18667), .n410(n410), .n18815(n18815), .n31(n31), 
            .n321(n321), .n6_adj_13(n6), .pwm_out2_c(pwm_out2_c), .\cycle_17__N_663[7] (cycle_17__N_663[7]), 
            .n14_adj_14(n14_adj_1471), .n3(n3_adj_1473), .\cycle_17__N_740[12] (cycle_17__N_740[12]), 
            .n18772(n18772), .n3_adj_15(n3), .\cycle_17__N_740[11] (cycle_17__N_740[11]), 
            .n7_adj_16(n7_adj_1472), .n18734(n18734), .\key_value[7] (key_value[7]), 
            .\key_value[9] (key_value[9]), .n18758(n18758), .\key_value[8] (key_value[8]), 
            .\key_flag[11] (key_flag[11]), .n18771(n18771), .n18814(n18814), 
            .n18768(n18768), .n18620(n18620), .n5_adj_17(n5), .\key_flag[12] (key_flag[12]), 
            .n18709(n18709), .n18770(n18770), .\key_value[0] (key_value[0]), 
            .n18685(n18685), .n18619(n18619), .n16876(n16876), .clk_N_168_enable_512(clk_N_168_enable_512), 
            .n18736(n18736), .n18735(n18735), .n18725(n18725), .n247(n247), 
            .n18708(n18708), .n9(n9), .n331(n331), .n415(n415), .n18651(n18651), 
            .n18308(n18308), .n18850(n18850), .\key_value[2] (key_value[2]), 
            .\key_value[3] (key_value[3]), .\key_value[6] (key_value[6]), 
            .n26_adj_18(n26_adj_1436), .\cycle_17__N_663[2] (cycle_17__N_663[2]), 
            .n10337(n10337), .n18707(n18707), .n269(n269), .n22_adj_19(n22_adj_1437), 
            .n18769(n18769), .n16920(n16920), .n18612(n18612), .n16959(n16959), 
            .n18623(n18623), .n417(n417), .\cycle_17__N_740[1] (cycle_17__N_740[1]), 
            .n18697(n18697), .\cycle_17__N_740[14] (cycle_17__N_740[14]), 
            .n19_adj_20(n19_adj_1438), .n17110(n17110), .n12983(n12983), 
            .n9757(n9757), .n17135(n17135), .\PWM_in_12__N_452[12] (PWM_in_12__N_452[12]), 
            .n37(n37), .n464(n464), .\key_flag[3] (key_flag[3]), .\key_flag[5] (key_flag[5]), 
            .\key_flag[6] (key_flag[6]), .n18756(n18756), .n34(n34), .en_1__N_194(en_1__N_194), 
            .n18606(n18606), .n18721(n18721), .n18668(n18668), .n3815(n3815), 
            .n3830(n3830), .n3800(n3800), .\key_flag[4] (key_flag[4]), 
            .\key_flag[7] (key_flag[7]), .n18684(n18684), .n18682(n18682), 
            .n16828(n16828), .n18706(n18706), .n16888(n16888), .n18616(n18616), 
            .\cycle_17__N_740[3] (cycle_17__N_740[3]), .n414(n414), .\cycle_17__N_740[4] (cycle_17__N_740[4]), 
            .\cycle_17__N_740[16] (cycle_17__N_740[16]), .n405(n405), .\cycle_17__N_740[13] (cycle_17__N_740[13]), 
            .n262(n262), .\cycle_17__N_740[9] (cycle_17__N_740[9]), .\PWM_in_12__N_452[10] (PWM_in_12__N_452[10]), 
            .\PWM_in_12__N_452[11] (PWM_in_12__N_452[11]), .\PWM_in_12__N_452[8] (PWM_in_12__N_452[8]), 
            .\PWM_in_12__N_452[9] (PWM_in_12__N_452[9]), .\PWM_in_12__N_452[6] (PWM_in_12__N_452[6]), 
            .\PWM_in_12__N_452[7] (PWM_in_12__N_452[7]), .\PWM_in_12__N_452[4] (PWM_in_12__N_452[4]), 
            .\PWM_in_12__N_452[5] (PWM_in_12__N_452[5]), .n58(n58), .n351(n351), 
            .n18655(n18655), .n18680(n18680), .clk_N_168_enable_507(clk_N_168_enable_507), 
            .clk_N_168_enable_518(clk_N_168_enable_518), .n17234(n17234), 
            .n17235(n17235), .n18785(n18785), .n18784(n18784), .n18757(n18757), 
            .n18717(n18717), .n19839(n19839), .\fcw_r_15__N_495[11] (fcw_r_15__N_495_adj_1733[11]), 
            .\fcw_r_15__N_495[5] (fcw_r_15__N_495_adj_1720[5]), .n8147(n8147), 
            .n8146(n8146), .yinjie({yinjie}), .clk__inv(clk__inv), .\fcw_r_15__N_495[9] (fcw_r_15__N_495_adj_1720[9]), 
            .clk(clk), .rst_n_c(rst_n_c), .key_pa_c(key_pa_c), .\fcw_r_15__N_495[10] (fcw_r_15__N_495_adj_1720[10]), 
            .\fcw_r_15__N_495[6] (fcw_r_15__N_495_adj_1720[6]), .\fcw_r_15__N_495[8] (fcw_r_15__N_495_adj_1720[8]), 
            .n18690(n18690), .n10972(n10972), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(36[9] 45[3])
    key u_key_state (.clk_N_168(clk_N_168), .key_state_flag(key_state_flag), 
        .key_state_c(key_state_c), .key_state_value(key_state_value), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(172[5] 178[4])
    IB key_pad_11 (.I(key[11]), .O(key_c_11));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    CCU2D cnt_2220_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15785), 
          .COUT(n15786), .S0(n128), .S1(n127));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_7.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_7.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_7.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_7.INJECT1_1 = "NO";
    IB key_pad_12 (.I(key[12]), .O(key_c_12));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_13 (.I(key[13]), .O(key_c_13));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_14 (.I(key[14]), .O(key_c_14));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // d:/fpga_project/lattice_diamond/piano/piano.v(4[9:14])
    IB sys_clk_pad (.I(sys_clk), .O(sys_clk_c));   // d:/fpga_project/lattice_diamond/piano/piano.v(3[12:19])
    OB pwm_out2_pad (.I(pwm_out2_c), .O(pwm_out2));   // d:/fpga_project/lattice_diamond/piano/piano.v(9[10:18])
    OB pwm_out1_pad (.I(pwm_out1_c), .O(pwm_out1));   // d:/fpga_project/lattice_diamond/piano/piano.v(8[10:18])
    CCU2D cnt_2220_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15784), 
          .COUT(n15785), .S0(n130), .S1(n129));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_5.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_5.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_5.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_5.INJECT1_1 = "NO";
    CCU2D cnt_2220_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15783), 
          .COUT(n15784), .S0(n132), .S1(n131));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_3.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_3.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_3.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_3.INJECT1_1 = "NO";
    CCU2D cnt_2220_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15783), .S1(n133));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_1.INIT0 = 16'hF000;
    defparam cnt_2220_add_4_1.INIT1 = 16'h0555;
    defparam cnt_2220_add_4_1.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_1.INJECT1_1 = "NO";
    LUT4 i7458_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n95), 
         .Z(n115)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7458_2_lut_3_lut.init = 16'hd0d0;
    CCU2D count_note_2222_add_4_9 (.A0(count_note[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15708), .S0(n38_adj_1457));   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222_add_4_9.INIT0 = 16'hfaaa;
    defparam count_note_2222_add_4_9.INIT1 = 16'h0000;
    defparam count_note_2222_add_4_9.INJECT1_0 = "NO";
    defparam count_note_2222_add_4_9.INJECT1_1 = "NO";
    CCU2D count_note_2222_add_4_7 (.A0(count_note[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_note[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15707), .COUT(n15708), .S0(n40_adj_1456), 
          .S1(n39));   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222_add_4_7.INIT0 = 16'hfaaa;
    defparam count_note_2222_add_4_7.INIT1 = 16'hfaaa;
    defparam count_note_2222_add_4_7.INJECT1_0 = "NO";
    defparam count_note_2222_add_4_7.INJECT1_1 = "NO";
    CCU2D count_note_2222_add_4_5 (.A0(count_note[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_note[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15706), .COUT(n15707), .S0(n42_adj_1454), 
          .S1(n41_adj_1455));   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222_add_4_5.INIT0 = 16'hfaaa;
    defparam count_note_2222_add_4_5.INIT1 = 16'hfaaa;
    defparam count_note_2222_add_4_5.INJECT1_0 = "NO";
    defparam count_note_2222_add_4_5.INJECT1_1 = "NO";
    CCU2D count_note_2222_add_4_3 (.A0(count_note[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_note[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15705), .COUT(n15706), .S0(n44_adj_1453), 
          .S1(n43));   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222_add_4_3.INIT0 = 16'hfaaa;
    defparam count_note_2222_add_4_3.INIT1 = 16'hfaaa;
    defparam count_note_2222_add_4_3.INJECT1_0 = "NO";
    defparam count_note_2222_add_4_3.INJECT1_1 = "NO";
    CCU2D count_note_2222_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_note[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n15705), .S1(n45));   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222_add_4_1.INIT0 = 16'hF000;
    defparam count_note_2222_add_4_1.INIT1 = 16'h0555;
    defparam count_note_2222_add_4_1.INJECT1_0 = "NO";
    defparam count_note_2222_add_4_1.INJECT1_1 = "NO";
    PFUMX i12620 (.BLUT(n18845), .ALUT(n18846), .C0(count_note[0]), .Z(n18847));
    LUT4 mux_617_Mux_0_i7_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[1]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n7_adj_1441)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !((C+!(D))+!B)) */ ;
    defparam mux_617_Mux_0_i7_4_lut_4_lut_4_lut.init = 16'hae02;
    LUT4 mux_617_Mux_2_i22_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n22_adj_1464)) /* synthesis lut_function=(A (B (D)+!B !(C+(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_617_Mux_2_i22_4_lut_4_lut_4_lut.init = 16'hdc07;
    LUT4 i11938_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[3]), 
         .C(count_note[0]), .D(count_note[1]), .Z(n17229)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (C+(D))+!B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11938_4_lut_4_lut_4_lut.init = 16'h5542;
    LUT4 i11849_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[3]), 
         .C(count_note[0]), .D(count_note[1]), .Z(n17140)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+!(D)))+!A (B+(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11849_4_lut_4_lut_4_lut.init = 16'hd65d;
    LUT4 mux_674_Mux_2_i7_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[3]), 
         .C(count_note[0]), .D(count_note[1]), .Z(n7)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_674_Mux_2_i7_4_lut_4_lut_4_lut.init = 16'h0540;
    L6MUX21 i12547 (.D0(n18461), .D1(n18458), .SD(count_note[4]), .Z(n18462));
    LUT4 i11861_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[3]), 
         .C(count_note[0]), .D(count_note[1]), .Z(n17152)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B+!(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11861_4_lut_4_lut_4_lut.init = 16'h6f64;
    LUT4 i12109_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n70_adj_1505)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i12109_3_lut_4_lut_4_lut_4_lut.init = 16'hfd7e;
    LUT4 count_note_5__bdd_4_lut_4_lut (.A(count_note[5]), .B(count_note[1]), 
         .C(count_note[0]), .D(count_note[2]), .Z(n18460)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A !(B+(C+(D))))) */ ;
    defparam count_note_5__bdd_4_lut_4_lut.init = 16'h7f76;
    LUT4 i12046_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[2]), 
         .C(count_note[1]), .D(count_note[3]), .Z(n17200)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C (D))+!B (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i12046_3_lut_4_lut_4_lut.init = 16'ha7f6;
    LUT4 i12065_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17151)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i12065_3_lut_4_lut_4_lut.init = 16'hb489;
    LUT4 i5564_3_lut_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n10407)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A !(B (C+(D))+!B ((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i5564_3_lut_3_lut_4_lut_4_lut.init = 16'h77e9;
    LUT4 mux_674_Mux_2_i14_3_lut_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), 
         .B(count_note[1]), .C(count_note[2]), .D(count_note[3]), .Z(n14_adj_1440)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B+!(C (D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam mux_674_Mux_2_i14_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1080;
    LUT4 mux_617_Mux_4_i92_3_lut_4_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n92_adj_1474)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_4_i92_3_lut_4_lut_4_lut_4_lut.init = 16'hc898;
    LUT4 mux_617_Mux_3_i7_3_lut_4_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n7_adj_1461)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_3_i7_3_lut_4_lut_4_lut_4_lut.init = 16'h8386;
    LUT4 mux_617_Mux_3_i92_3_lut_3_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n92)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B (C (D))+!B !(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_3_i92_3_lut_3_lut_4_lut_4_lut.init = 16'h3477;
    LUT4 i10433_2_lut_rep_423_3_lut_4_lut (.A(n18760), .B(n18615), .C(n8_adj_1478), 
         .D(n18614), .Z(n18605)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i10433_2_lut_rep_423_3_lut_4_lut.init = 16'h8000;
    LUT4 i11932_4_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17223)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11932_4_lut_4_lut_4_lut_4_lut.init = 16'h6631;
    LUT4 i11903_3_lut_4_lut_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[1]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n17194)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A !((C+!(D))+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i11903_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h7bdd;
    LUT4 i11908_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17199)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C (D)+!C !(D))+!B (C+(D)))) */ ;
    defparam i11908_3_lut_4_lut_4_lut_4_lut.init = 16'hf1bc;
    LUT4 mux_617_Mux_3_i77_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n77_adj_1504)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_617_Mux_3_i77_3_lut_4_lut_4_lut_4_lut.init = 16'hf1a3;
    LUT4 mux_674_Mux_2_i29_3_lut_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), 
         .B(count_note[2]), .C(count_note[1]), .D(count_note[3]), .Z(n29)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((C+!(D))+!B))) */ ;
    defparam mux_674_Mux_2_i29_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0420;
    LUT4 mux_617_Mux_4_i22_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[2]), 
         .C(count_note[1]), .D(count_note[3]), .Z(n22_adj_1484)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)))+!A !(B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_617_Mux_4_i22_3_lut_4_lut_4_lut.init = 16'h83fb;
    LUT4 mux_617_Mux_1_i53_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n53)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C (D)+!C !(D))+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_1_i53_3_lut_4_lut_4_lut.init = 16'h0442;
    PFUMX i12542 (.BLUT(n17173), .ALUT(n18457), .C0(count_note[5]), .Z(n18458));
    LUT4 i29_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[4]), .Z(n16_adj_1439)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i29_3_lut_4_lut_4_lut.init = 16'h04c7;
    CCU2D sub_1378_add_2_19 (.A0(CNT[17]), .B0(CNT_17__N_703[17]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15507), .S1(n3759));
    defparam sub_1378_add_2_19.INIT0 = 16'h5999;
    defparam sub_1378_add_2_19.INIT1 = 16'h0000;
    defparam sub_1378_add_2_19.INJECT1_0 = "NO";
    defparam sub_1378_add_2_19.INJECT1_1 = "NO";
    LUT4 mux_674_Mux_1_i7_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n7_adj_1503)) /* synthesis lut_function=(A (B+(C+!(D)))+!A ((C)+!B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam mux_674_Mux_1_i7_4_lut_4_lut.init = 16'hf9fb;
    CCU2D sub_1378_add_2_17 (.A0(CNT[15]), .B0(CNT_17__N_703[15]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[16]), .B1(CNT_17__N_703[16]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15506), .COUT(n15507));
    defparam sub_1378_add_2_17.INIT0 = 16'h5999;
    defparam sub_1378_add_2_17.INIT1 = 16'h5999;
    defparam sub_1378_add_2_17.INJECT1_0 = "NO";
    defparam sub_1378_add_2_17.INJECT1_1 = "NO";
    LUT4 mux_617_Mux_2_i14_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n14_adj_1466)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_2_i14_3_lut_4_lut.init = 16'h983d;
    LUT4 mux_617_Mux_0_i101_3_lut_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n101_adj_1511)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(B (C+(D))+!B (C (D)))) */ ;
    defparam mux_617_Mux_0_i101_3_lut_3_lut_4_lut_4_lut.init = 16'ha31f;
    LUT4 mux_617_Mux_4_i7_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n7_adj_1486)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam mux_617_Mux_4_i7_3_lut_4_lut_4_lut.init = 16'h3de0;
    CCU2D sub_1378_add_2_15 (.A0(CNT[13]), .B0(CNT_17__N_703[13]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[14]), .B1(CNT_17__N_703[14]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15505), .COUT(n15506));
    defparam sub_1378_add_2_15.INIT0 = 16'h5999;
    defparam sub_1378_add_2_15.INIT1 = 16'h5999;
    defparam sub_1378_add_2_15.INJECT1_0 = "NO";
    defparam sub_1378_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_1378_add_2_13 (.A0(CNT[11]), .B0(CNT_17__N_703[11]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[12]), .B1(CNT_17__N_703[12]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15504), .COUT(n15505));
    defparam sub_1378_add_2_13.INIT0 = 16'h5999;
    defparam sub_1378_add_2_13.INIT1 = 16'h5999;
    defparam sub_1378_add_2_13.INJECT1_0 = "NO";
    defparam sub_1378_add_2_13.INJECT1_1 = "NO";
    LUT4 mux_617_Mux_0_i70_3_lut_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n70)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C))) */ ;
    defparam mux_617_Mux_0_i70_3_lut_3_lut_4_lut_4_lut.init = 16'h9d1f;
    LUT4 i11910_3_lut (.A(n37_adj_1467), .B(n91), .C(count_note[3]), .Z(n17201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11910_3_lut.init = 16'hcaca;
    LUT4 i11850_4_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n17141)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i11850_4_lut_4_lut_4_lut.init = 16'h27b0;
    LUT4 mux_617_Mux_0_i77_3_lut_4_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n77)) /* synthesis lut_function=(A ((C)+!B)+!A (B+((D)+!C))) */ ;
    defparam mux_617_Mux_0_i77_3_lut_4_lut_4_lut_4_lut.init = 16'hf7e7;
    LUT4 n17173_bdd_4_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n18457)) /* synthesis lut_function=(!(A (B+(C))+!A (B (C)+!B !((D)+!C)))) */ ;
    defparam n17173_bdd_4_lut_4_lut_4_lut.init = 16'h1707;
    LUT4 i7946_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n83), 
         .Z(n103)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7946_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_617_Mux_0_i92_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n92_adj_1512)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B (C)+!B !(C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_0_i92_3_lut_4_lut_4_lut.init = 16'he3f9;
    LUT4 mux_617_Mux_3_i38_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n38_adj_1462)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A (B+!(C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_3_i38_3_lut_4_lut_4_lut.init = 16'hcf7d;
    PFUMX i12545 (.BLUT(n18460), .ALUT(n18459), .C0(count_note[3]), .Z(n18461));
    LUT4 i11876_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17167)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A !(D))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11876_4_lut_4_lut_4_lut.init = 16'h7da8;
    CCU2D sub_1378_add_2_11 (.A0(CNT[9]), .B0(CNT_17__N_703[9]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[10]), .B1(CNT_17__N_703[10]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15503), .COUT(n15504));
    defparam sub_1378_add_2_11.INIT0 = 16'h5999;
    defparam sub_1378_add_2_11.INIT1 = 16'h5999;
    defparam sub_1378_add_2_11.INJECT1_0 = "NO";
    defparam sub_1378_add_2_11.INJECT1_1 = "NO";
    LUT4 mux_617_Mux_3_i53_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n53_adj_1508)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+!(D)))+!A !(B (C+(D))+!B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_3_i53_3_lut_4_lut_4_lut.init = 16'h7de2;
    LUT4 i11848_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n17139)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C))) */ ;
    defparam i11848_3_lut_4_lut.init = 16'he94d;
    CCU2D sub_1378_add_2_9 (.A0(CNT[7]), .B0(CNT_17__N_703[7]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[8]), .B1(CNT_17__N_703[8]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15502), .COUT(n15503));
    defparam sub_1378_add_2_9.INIT0 = 16'h5999;
    defparam sub_1378_add_2_9.INIT1 = 16'h5999;
    defparam sub_1378_add_2_9.INJECT1_0 = "NO";
    defparam sub_1378_add_2_9.INJECT1_1 = "NO";
    LUT4 i12067_3_lut_4_lut (.A(count_note[2]), .B(count_note[1]), .C(count_note[0]), 
         .D(count_note[3]), .Z(n17149)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i12067_3_lut_4_lut.init = 16'h4974;
    CCU2D sub_1378_add_2_7 (.A0(CNT[5]), .B0(CNT_17__N_703[5]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[6]), .B1(CNT_17__N_703[6]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15501), .COUT(n15502));
    defparam sub_1378_add_2_7.INIT0 = 16'h5999;
    defparam sub_1378_add_2_7.INIT1 = 16'h5999;
    defparam sub_1378_add_2_7.INJECT1_0 = "NO";
    defparam sub_1378_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_1378_add_2_5 (.A0(CNT[3]), .B0(CNT_17__N_703[3]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[4]), .B1(CNT_17__N_703[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15500), .COUT(n15501));
    defparam sub_1378_add_2_5.INIT0 = 16'h5999;
    defparam sub_1378_add_2_5.INIT1 = 16'h5999;
    defparam sub_1378_add_2_5.INJECT1_0 = "NO";
    defparam sub_1378_add_2_5.INJECT1_1 = "NO";
    FD1S3AX count_beat_i4_2224__i0 (.D(n30_adj_1481), .CK(clk_N_168), .Q(count_beat[0]));   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam count_beat_i4_2224__i0.GSR = "DISABLED";
    LUT4 mux_674_Mux_1_i29_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n29_adj_1458)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_674_Mux_1_i29_4_lut_4_lut_4_lut.init = 16'hebf7;
    LUT4 mux_617_Mux_4_i45_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n45_adj_1482)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A !(B+(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_4_i45_3_lut_4_lut_4_lut.init = 16'h8102;
    LUT4 i11859_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17150)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11859_3_lut_4_lut_4_lut.init = 16'h7a4b;
    LUT4 i11851_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17142)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(B (C)+!B !(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11851_3_lut_4_lut_4_lut.init = 16'h4be9;
    LUT4 i11875_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17166)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11875_3_lut_4_lut_4_lut.init = 16'hfe69;
    LUT4 i7941_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n88), 
         .Z(n108)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7941_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i11874_3_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[0]), 
         .C(count_note[1]), .D(count_note[3]), .Z(n17165)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A ((C)+!B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11874_3_lut_4_lut_4_lut.init = 16'hf17b;
    LUT4 i11877_3_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[0]), 
         .C(count_note[1]), .D(count_note[3]), .Z(n17168)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11877_3_lut_4_lut_4_lut.init = 16'h69f1;
    CCU2D sub_1378_add_2_3 (.A0(CNT[1]), .B0(CNT_17__N_703[1]), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[2]), .B1(CNT_17__N_703[2]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15499), .COUT(n15500));
    defparam sub_1378_add_2_3.INIT0 = 16'h5999;
    defparam sub_1378_add_2_3.INIT1 = 16'h5999;
    defparam sub_1378_add_2_3.INJECT1_0 = "NO";
    defparam sub_1378_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_1378_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[0]), .B1(CNT_17__N_703[0]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15499));
    defparam sub_1378_add_2_1.INIT0 = 16'h0000;
    defparam sub_1378_add_2_1.INIT1 = 16'h5999;
    defparam sub_1378_add_2_1.INJECT1_0 = "NO";
    defparam sub_1378_add_2_1.INJECT1_1 = "NO";
    LUT4 i11901_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17192)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i11901_3_lut_4_lut_4_lut.init = 16'hae7b;
    LUT4 i11907_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17198)) /* synthesis lut_function=(!(A (B (D))+!A !(B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam i11907_3_lut_4_lut_4_lut.init = 16'h67ae;
    LUT4 i11930_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17221)) /* synthesis lut_function=(A (B (D))+!A !(B ((D)+!C)+!B !(C+!(D)))) */ ;
    defparam i11930_3_lut_4_lut_4_lut.init = 16'h9851;
    LUT4 i11902_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n17193)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i11902_3_lut_4_lut.init = 16'h79e4;
    LUT4 i11922_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n17213)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A (B (D)+!B !(D))) */ ;
    defparam i11922_3_lut_4_lut.init = 16'hc61b;
    LUT4 i11931_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n17222)) /* synthesis lut_function=(A (B (D)+!B !(C (D)))+!A !(B (C (D)+!C !(D))+!B (C+(D)))) */ ;
    defparam i11931_3_lut_4_lut.init = 16'h8e63;
    LUT4 i11937_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n17228)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B+!(C (D)+!C !(D))))) */ ;
    defparam i11937_3_lut_4_lut.init = 16'h1a81;
    LUT4 i12037_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n17224)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B (D)+!B !(D))) */ ;
    defparam i12037_3_lut_4_lut.init = 16'he639;
    FD1P3AX stat_71 (.D(n17430), .SP(VCC_net), .CK(clk__inv), .Q(stat)) /* synthesis lse_init_val=0 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(196[7] 205[5])
    defparam stat_71.GSR = "ENABLED";
    LUT4 i7947_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n82), 
         .Z(n102)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7947_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7948_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n81), 
         .Z(n101)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7948_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7937_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n92_adj_1476), 
         .Z(n112)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7937_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7949_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n80), 
         .Z(n100)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7949_2_lut_3_lut.init = 16'hd0d0;
    PFUMX i12536 (.BLUT(n18442), .ALUT(n18441), .C0(count_note[5]), .Z(n18443));
    LUT4 LessThan_51_i4_4_lut (.A(beat[0]), .B(beat[1]), .C(count_beat[1]), 
         .D(count_beat[0]), .Z(n4_adj_1452)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(242[8:25])
    defparam LessThan_51_i4_4_lut.init = 16'h0c8e;
    LUT4 i2331_3_lut_rep_487 (.A(yinjie[0]), .B(n73), .C(n10074), .Z(n18669)) /* synthesis lut_function=(A+!(B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(213[7] 218[5])
    defparam i2331_3_lut_rep_487.init = 16'habab;
    LUT4 i1_3_lut_4_lut (.A(yinjie[0]), .B(n73), .C(n10074), .D(yinjie[1]), 
         .Z(n13)) /* synthesis lut_function=(A ((D)+!B)+!A !(B+!((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(213[7] 218[5])
    defparam i1_3_lut_4_lut.init = 16'hbb23;
    FD1S3IX cnt_2220__i0 (.D(n133), .CK(clk_N_168), .CD(n10969), .Q(cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i0.GSR = "ENABLED";
    LUT4 i2_4_lut_4_lut (.A(n73), .B(n19846), .C(yinjie[1]), .D(n18669), 
         .Z(yinjie_2__N_1[1])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam i2_4_lut_4_lut.init = 16'hd2e1;
    LUT4 i2_4_lut_4_lut_adj_56 (.A(n73), .B(n19846), .C(yinjie[2]), .D(n13), 
         .Z(yinjie_2__N_1[2])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam i2_4_lut_4_lut_adj_56.init = 16'hd2e1;
    LUT4 i1_4_lut (.A(n41), .B(cnt[15]), .C(n46), .D(n42), .Z(n9_adj_1506)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i11716_4_lut (.A(cnt[13]), .B(cnt[9]), .C(cnt[22]), .D(cnt[11]), 
         .Z(n17005)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11716_4_lut.init = 16'h8000;
    LUT4 i17_4_lut (.A(cnt[24]), .B(cnt[19]), .C(cnt[16]), .D(cnt[21]), 
         .Z(n41)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(n25_adj_1450), .B(n44), .C(n38), .D(n26_adj_1449), 
         .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(cnt[26]), .B(cnt[8]), .C(cnt[10]), .D(cnt[14]), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i18_4_lut.init = 16'hfffe;
    FD1P3IX count_note_2222__i0 (.D(n45), .SP(clk_N_168_enable_533), .CD(n10968), 
            .CK(clk_N_168), .Q(count_note[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i0.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(cnt[7]), .B(cnt[4]), .Z(n25_adj_1450)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i20_4_lut (.A(cnt[2]), .B(n40), .C(n30), .D(cnt[31]), .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(cnt[30]), .B(cnt[20]), .C(cnt[6]), .D(cnt[1]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i7950_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n79), 
         .Z(n99)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7950_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i2_2_lut (.A(cnt[23]), .B(cnt[29]), .Z(n26_adj_1449)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i7951_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n78), 
         .Z(n98)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7951_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i8154_3_lut_3_lut (.A(count_note[3]), .B(count_note[1]), .C(count_note[2]), 
         .Z(n13008)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam i8154_3_lut_3_lut.init = 16'hd0d0;
    LUT4 i16_4_lut (.A(cnt[28]), .B(cnt[12]), .C(cnt[3]), .D(cnt[17]), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(cnt[27]), .B(cnt[25]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i12325_4_lut (.A(n18812), .B(n16847), .C(count_note[5]), .D(count_note[4]), 
         .Z(clk_N_168_enable_456)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam i12325_4_lut.init = 16'h373f;
    FD1P3AX beat_i2 (.D(beat_4__N_40[2]), .SP(clk_N_168_enable_456), .CK(clk_N_168), 
            .Q(beat[2]));   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam beat_i2.GSR = "DISABLED";
    FD1P3AX beat_i1 (.D(beat_4__N_40[1]), .SP(clk_N_168_enable_456), .CK(clk_N_168), 
            .Q(beat[1]));   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam beat_i1.GSR = "DISABLED";
    FD1P3AX note_i4 (.D(note_5__N_45[4]), .SP(clk_N_168_enable_534), .CK(clk_N_168), 
            .Q(note[4]));   // d:/fpga_project/lattice_diamond/piano/piano.v(255[7] 514[4])
    defparam note_i4.GSR = "DISABLED";
    FD1P3AX note_i3 (.D(note_5__N_45[3]), .SP(clk_N_168_enable_534), .CK(clk_N_168), 
            .Q(note[3]));   // d:/fpga_project/lattice_diamond/piano/piano.v(255[7] 514[4])
    defparam note_i3.GSR = "DISABLED";
    FD1P3AX note_i2 (.D(note_5__N_45[2]), .SP(clk_N_168_enable_456), .CK(clk_N_168), 
            .Q(note[2]));   // d:/fpga_project/lattice_diamond/piano/piano.v(255[7] 514[4])
    defparam note_i2.GSR = "DISABLED";
    FD1P3AX note_i1 (.D(note_5__N_45[1]), .SP(clk_N_168_enable_456), .CK(clk_N_168), 
            .Q(note[1]));   // d:/fpga_project/lattice_diamond/piano/piano.v(255[7] 514[4])
    defparam note_i1.GSR = "DISABLED";
    LUT4 i11919_3_lut (.A(n17208), .B(n17209), .C(count_note[7]), .Z(note_5__N_45[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11919_3_lut.init = 16'hcaca;
    LUT4 i11918_3_lut (.A(n17148), .B(n109_adj_1509), .C(count_note[6]), 
         .Z(n17209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11918_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_57 (.A(count_note[7]), .B(count_note[6]), .Z(n16847)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_57.init = 16'h8888;
    LUT4 i12370_3_lut_2_lut_3_lut (.A(key_state_flag), .B(key_state_value), 
         .C(n19846), .Z(n17430)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(198[7:41])
    defparam i12370_3_lut_2_lut_3_lut.init = 16'hd2d2;
    LUT4 i2_4_lut (.A(n73), .B(n10074), .C(n19846), .D(yinjie[0]), .Z(yinjie_2__N_1[0])) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i2_4_lut.init = 16'hf10e;
    LUT4 i3_4_lut (.A(key_value[14]), .B(n12259), .C(key_flag[14]), .D(yinjie[2]), 
         .Z(n73)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i11711_3_lut_4_lut (.A(count_note[3]), .B(n18779), .C(count_note[4]), 
         .D(count_note[5]), .Z(n6_adj_1488)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i11711_3_lut_4_lut.init = 16'h0002;
    LUT4 i12338_4_lut (.A(count_note[5]), .B(n16847), .C(n18671), .D(count_note[4]), 
         .Z(clk_N_168_enable_534)) /* synthesis lut_function=(!(A (B)+!A (B (C (D))))) */ ;
    defparam i12338_4_lut.init = 16'h3777;
    LUT4 i2_4_lut_adj_58 (.A(n16854), .B(count_note[0]), .C(n18604), .D(count_note[4]), 
         .Z(beat_4__N_40[4])) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i2_4_lut_adj_58.init = 16'h3200;
    LUT4 i7940_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n89), 
         .Z(n109)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7940_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i683_2_lut_rep_578 (.A(clk_beat), .B(n19846), .Z(n18760)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(240[3] 252[9])
    defparam i683_2_lut_rep_578.init = 16'h8888;
    LUT4 i10415_2_lut_3_lut_4_lut (.A(clk_beat), .B(n19846), .C(n4689), 
         .D(count_beat[0]), .Z(n30_adj_1481)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(240[3] 252[9])
    defparam i10415_2_lut_3_lut_4_lut.init = 16'h7888;
    LUT4 i10417_2_lut_rep_425_3_lut_4_lut (.A(clk_beat), .B(n19846), .C(n4689), 
         .D(count_beat[0]), .Z(n18607)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(240[3] 252[9])
    defparam i10417_2_lut_rep_425_3_lut_4_lut.init = 16'h8000;
    LUT4 i2098_2_lut_3_lut (.A(clk_beat), .B(n19846), .C(n201), .Z(n4689)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(240[3] 252[9])
    defparam i2098_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i10437_2_lut_3_lut_4_lut (.A(n18614), .B(n18607), .C(n18613), 
         .D(n8_adj_1478), .Z(n27)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i10437_2_lut_3_lut_4_lut.init = 16'h78f0;
    IB key_pad_8 (.I(key[8]), .O(key_c_8));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_7 (.I(key[7]), .O(key_c_7));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_6 (.I(key[6]), .O(key_c_6));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_5 (.I(key[5]), .O(key_c_5));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_4 (.I(key[4]), .O(key_c_4));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_3 (.I(key[3]), .O(key_c_3));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_2 (.I(key[2]), .O(key_c_2));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_1 (.I(key[1]), .O(key_c_1));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pad_0 (.I(key[0]), .O(key_c_0));   // d:/fpga_project/lattice_diamond/piano/piano.v(5[16:19])
    IB key_pa_pad (.I(key_pa), .O(key_pa_c));   // d:/fpga_project/lattice_diamond/piano/piano.v(6[9:15])
    IB key_state_pad (.I(key_state), .O(key_state_c));   // d:/fpga_project/lattice_diamond/piano/piano.v(7[9:18])
    LUT4 mux_617_Mux_1_i38_3_lut_4_lut (.A(count_note[0]), .B(n18773), .C(count_note[3]), 
         .D(n37_adj_1467), .Z(n38_adj_1468)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_1_i38_3_lut_4_lut.init = 16'hf404;
    PFUMX i12618 (.BLUT(n18842), .ALUT(n18843), .C0(count_note[0]), .Z(n18844));
    LUT4 i7954_2_lut_rep_431 (.A(count_beat[3]), .B(n4689), .Z(n18613)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i7954_2_lut_rep_431.init = 16'h8888;
    PFUMX i12616 (.BLUT(n18839), .ALUT(n18840), .C0(count_note[0]), .Z(n18841));
    LUT4 i1_2_lut_rep_591 (.A(count_note[1]), .B(count_note[2]), .Z(n18773)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i1_2_lut_rep_591.init = 16'h2222;
    LUT4 i2_2_lut_3_lut (.A(count_note[1]), .B(count_note[2]), .C(count_note[3]), 
         .Z(n7_adj_1448)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i2_2_lut_3_lut.init = 16'h2020;
    LUT4 count_note_5__bdd_2_lut_12560_3_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[4]), .Z(n18441)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam count_note_5__bdd_2_lut_12560_3_lut.init = 16'h0202;
    LUT4 i8169_3_lut_4_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n13024)) /* synthesis lut_function=(!(A (B (C)+!B !(C+!(D)))+!A (B (C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i8169_3_lut_4_lut_4_lut.init = 16'h3d3f;
    LUT4 i1_2_lut_rep_592 (.A(count_note[0]), .B(count_note[3]), .Z(n18774)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_592.init = 16'hbbbb;
    LUT4 i2_3_lut_3_lut_4_lut (.A(count_note[0]), .B(count_note[3]), .C(count_note[2]), 
         .D(count_note[1]), .Z(n16896)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i2_3_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 i8113_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[3]), 
         .D(count_note[2]), .Z(n45_adj_1469)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;
    defparam i8113_3_lut_4_lut.init = 16'h1001;
    LUT4 i1_2_lut_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[3]), 
         .D(count_note[2]), .Z(n16860)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i5562_3_lut_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n10405)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A (B+!((D)+!C)))) */ ;
    defparam i5562_3_lut_3_lut_4_lut.init = 16'h33a1;
    LUT4 i10444_4_lut_4_lut (.A(count_beat[3]), .B(n4689), .C(n18605), 
         .D(count_beat[4]), .Z(n26_adj_1479)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A !(B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i10444_4_lut_4_lut.init = 16'h4c80;
    LUT4 i7407_2_lut (.A(yinjie[0]), .B(yinjie[1]), .Z(n12259)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7407_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_597 (.A(count_note[2]), .B(count_note[1]), .Z(n18779)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i1_2_lut_rep_597.init = 16'hdddd;
    LUT4 count_note_5__bdd_3_lut_12544_4_lut (.A(count_note[2]), .B(count_note[1]), 
         .C(count_note[4]), .D(count_note[0]), .Z(n18442)) /* synthesis lut_function=(!((B+!(C (D)+!C !(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam count_note_5__bdd_3_lut_12544_4_lut.init = 16'h2002;
    LUT4 i2_4_lut_adj_59 (.A(yinjie[1]), .B(key_value[13]), .C(yinjie[2]), 
         .D(key_flag[13]), .Z(n10074)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(214[6:55])
    defparam i2_4_lut_adj_59.init = 16'h3200;
    LUT4 i7952_2_lut_rep_432 (.A(count_beat[1]), .B(n4689), .Z(n18614)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i7952_2_lut_rep_432.init = 16'h8888;
    LUT4 i7468_3_lut_3_lut_4_lut (.A(count_note[2]), .B(count_note[1]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n10403)) /* synthesis lut_function=(!((B+!(C (D)+!C !(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i7468_3_lut_3_lut_4_lut.init = 16'h2002;
    LUT4 count_note_5__bdd_3_lut_12551_4_lut (.A(count_note[2]), .B(count_note[1]), 
         .C(count_note[0]), .D(count_note[5]), .Z(n18459)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (C+!(D))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam count_note_5__bdd_3_lut_12551_4_lut.init = 16'hf2df;
    LUT4 i8026_2_lut_3_lut_4_lut (.A(count_note[2]), .B(count_note[1]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n38_adj_1483)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i8026_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_60 (.A(count_note[0]), .B(count_note[1]), .C(count_note[3]), 
         .D(count_note[2]), .Z(n16865)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_60.init = 16'h0220;
    LUT4 mux_617_Mux_1_i37_3_lut_3_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .Z(n37_adj_1467)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B (C))) */ ;
    defparam mux_617_Mux_1_i37_3_lut_3_lut.init = 16'hc2c2;
    LUT4 i12258_2_lut_rep_599 (.A(count_note[0]), .B(count_note[1]), .Z(n18781)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i12258_2_lut_rep_599.init = 16'h9999;
    LUT4 mux_674_Mux_1_i91_3_lut_3_lut_4_lut_3_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .Z(n91)) /* synthesis lut_function=(!(A (C)+!A (B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_674_Mux_1_i91_3_lut_3_lut_4_lut_3_lut.init = 16'h1b1b;
    LUT4 i1_2_lut_3_lut_4_lut_adj_61 (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n16868)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i1_2_lut_3_lut_4_lut_adj_61.init = 16'h000d;
    LUT4 i7938_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n91_adj_1475), 
         .Z(n111)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7938_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_617_Mux_0_i14_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n14)) /* synthesis lut_function=(A (B (D))+!A !(B (C)+!B !((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_0_i14_3_lut_4_lut_4_lut.init = 16'h9d05;
    LUT4 n18439_bdd_3_lut_then_4_lut (.A(count_note[5]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[4]), .Z(n18836)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B+!(C+!(D))))) */ ;
    defparam n18439_bdd_3_lut_then_4_lut.init = 16'h1231;
    LUT4 n18439_bdd_3_lut_else_4_lut (.A(count_note[5]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[4]), .Z(n18835)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(C (D)+!C !(D)))) */ ;
    defparam n18439_bdd_3_lut_else_4_lut.init = 16'h5085;
    LUT4 mux_617_Mux_0_i22_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n22_adj_1444)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B (C+(D))+!B (C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_0_i22_3_lut_4_lut_4_lut_4_lut.init = 16'h56f0;
    LUT4 i11920_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17211)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !(C (D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11920_3_lut_4_lut_4_lut_4_lut.init = 16'h30c6;
    LUT4 i7_4_lut (.A(n9_adj_1506), .B(n17005), .C(cnt[5]), .D(cnt[18]), 
         .Z(n10216)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i7_4_lut.init = 16'hbfff;
    buzzer u_buzzer (.CNT({CNT}), .GND_net(GND_net), .CNT_17__N_703({CNT_17__N_703}), 
           .clk_N_168(clk_N_168), .stat(stat), .\yinjie_box_2__N_394[0] (yinjie_box_2__N_394[0]), 
           .\yinjie_box_2__N_394[1] (yinjie_box_2__N_394[1]), .n77({n78, 
           n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
           n89, n90, n91_adj_1475, n92_adj_1476, n93, n94_adj_1477, 
           n95}), .n9292(n9292), .n19846(n19846), .\data_out2[0] (data_out2[0]), 
           .\data_out1[0] (data_out1[0]), .n28({n14_adj_1435, n15, n16, 
           n17, n18, n19, n20, n21, n22, n23, n24, n25, n26}), 
           .yinjie({yinjie}), .pwm_out1_c(pwm_out1_c), .\PWM_in_12__N_452[12] (PWM_in_12__N_452[12]), 
           .\PWM_in_12__N_452[11] (PWM_in_12__N_452[11]), .\PWM_in_12__N_452[10] (PWM_in_12__N_452[10]), 
           .\rom2[0] (rom2[0]), .n18850(n18850), .\PWM_in_12__N_452[9] (PWM_in_12__N_452[9]), 
           .n97({n98, n99, n100, n101, n102, n103, n104, n105, 
           n106, n107, n108, n109, n110, n111, n112, n113, n114, 
           n115}), .n18725(n18725), .n18707(n18707), .n18706(n18706), 
           .n18709(n18709), .n18721(n18721), .n18616(n18616), .\cycle_17__N_740[4] (cycle_17__N_740[4]), 
           .n17110(n17110), .n18755(n18755), .n18708(n18708), .n18736(n18736), 
           .n18684(n18684), .n7(n7_adj_1472), .\cycle_17__N_740[13] (cycle_17__N_740[13]), 
           .\PWM_in_12__N_452[8] (PWM_in_12__N_452[8]), .n407(n407), .\cycle_17__N_740[11] (cycle_17__N_740[11]), 
           .n18722(n18722), .n18763(n18763), .\cycle_17__N_740[14] (cycle_17__N_740[14]), 
           .n415(n415), .\cycle_17__N_740[3] (cycle_17__N_740[3]), .\note[0] (note[0]), 
           .n18737(n18737), .n18807(n18807), .n18697(n18697), .n18757(n18757), 
           .n18784(n18784), .n18785(n18785), .\fcw_r_15__N_495[8] (fcw_r_15__N_495_adj_1720[8]), 
           .\PWM_in_12__N_452[7] (PWM_in_12__N_452[7]), .n18690(n18690), 
           .\fcw_r_15__N_495[6] (fcw_r_15__N_495_adj_1720[6]), .n8146(n8146), 
           .n8147(n8147), .\fcw_r_15__N_495[10] (fcw_r_15__N_495_adj_1720[10]), 
           .\fcw_r_15__N_495[5] (fcw_r_15__N_495_adj_1720[5]), .n18717(n18717), 
           .n10972(n10972), .\fcw_r_15__N_495[11] (fcw_r_15__N_495_adj_1733[11]), 
           .\fcw_r_15__N_495[9] (fcw_r_15__N_495_adj_1720[9]), .n18620(n18620), 
           .n18668(n18668), .n16876(n16876), .\cycle_17__N_740[1] (cycle_17__N_740[1]), 
           .\note[1] (note[1]), .n18808(n18808), .n12983(n12983), .\PWM_in_12__N_452[6] (PWM_in_12__N_452[6]), 
           .\PWM_in_12__N_452[5] (PWM_in_12__N_452[5]), .n406(n406), .\cycle_17__N_740[12] (cycle_17__N_740[12]), 
           .clk_N_168_enable_507(clk_N_168_enable_507), .\cycle_17__N_663[2] (cycle_17__N_663[2]), 
           .clk_N_168_enable_512(clk_N_168_enable_512), .\cycle_17__N_663[7] (cycle_17__N_663[7]), 
           .\cycle_17__N_663[10] (cycle_17__N_663[10]), .clk_N_168_enable_518(clk_N_168_enable_518), 
           .\cycle_17__N_663[17] (cycle_17__N_663[17]), .\cycle_17__N_740[9] (cycle_17__N_740[9]), 
           .n18769(n18769), .\PWM_in_12__N_452[4] (PWM_in_12__N_452[4]), 
           .n19_adj_4(n19_adj_1438), .n22_adj_5(n22_adj_1437), .n18772(n18772), 
           .n14_adj_6(n14_adj_1471), .n3(n3), .n3_adj_7(n3_adj_1473), 
           .n18735(n18735), .n16828(n16828), .n18754(n18754), .n262(n262), 
           .\PWM_in_12__N_452[3] (PWM_in_12__N_452[3]), .n7_adj_8(n7_adj_1470), 
           .\cycle_17__N_740[16] (cycle_17__N_740[16]), .\PWM_in_12__N_452[2] (PWM_in_12__N_452[2]), 
           .n18720(n18720), .n18815(n18815), .n18651(n18651), .\PWM_in_12__N_452[1] (PWM_in_12__N_452[1]), 
           .n18803(n18803), .n18761(n18761), .n18768(n18768), .n18771(n18771), 
           .n18619(n18619), .clk__inv(clk__inv), .n410(n410), .n18623(n18623), 
           .\key_value[0] (key_value[0]), .\key_value[10] (key_value[10]), 
           .n269(n269), .n16959(n16959), .n26_adj_9(n26_adj_1436), .n9757(n9757), 
           .\cycle_17__N_740[10] (cycle_17__N_740[10]), .n18308(n18308), 
           .n18307(n18307), .\key_value[12] (key_value[12]), .\key_value[5] (key_value[5]), 
           .\key_value[1] (key_value[1]), .\key_value[8] (key_value[8]), 
           .\key_value[7] (key_value[7]), .\key_value[6] (key_value[6]), 
           .\key_value[2] (key_value[2]), .\key_value[11] (key_value[11]), 
           .\key_value[3] (key_value[3]), .\key_value[4] (key_value[4]), 
           .\key_value[9] (key_value[9]), .n3830(n3830), .n18679(n18679), 
           .n436(n436), .n18676(n18676), .\rom1_4__N_338[0] (rom1_4__N_338[0]), 
           .n351(n351), .n414(n414), .n31(n31), .n18682(n18682), .n16888(n16888), 
           .n18610(n18610), .n247(n247), .n331(n331), .\rom2[1] (rom2[1]), 
           .\key_flag[2] (key_flag[2]), .\key_flag[1] (key_flag[1]), .n18734(n18734), 
           .rst_n_c(rst_n_c), .key_pa_c(key_pa_c), .n19839(n19839), .n18680(n18680), 
           .n9(n9), .n9654(n9654), .n10160(n10160), .n344(n344), .n18696(n18696), 
           .n18606(n18606), .n18612(n18612), .n16920(n16920), .n10337(n10337), 
           .n18649(n18649), .n18685(n18685), .n18652(n18652), .n16909(n16909)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(182[8] 191[3])
    PFUMX i12614 (.BLUT(n18835), .ALUT(n18836), .C0(count_note[0]), .Z(n18837));
    L6MUX21 i11958 (.D0(n17164), .D1(n17171), .SD(count_note[6]), .Z(n17249));
    L6MUX21 i11917 (.D0(n17138), .D1(n17145), .SD(count_note[6]), .Z(n17208));
    L6MUX21 i11832 (.D0(n17207), .D1(n17217), .SD(count_note[6]), .Z(n17123));
    key_U17 u_key_5 (.clk_N_168(clk_N_168), .\key_flag[4] (key_flag[4]), 
            .key_c_4(key_c_4), .\key_value[4] (key_value[4]), .GND_net(GND_net), 
            .n18735(n18735), .n6(n6_adj_1443), .n5(n5_adj_1447), .n891(n891), 
            .n19846(n19846), .n18754(n18754), .n16888(n16888), .n18747(n18747), 
            .n5_adj_3(n5), .n11464(n11464), .n18722(n18722), .n18654(n18654), 
            .n18736(n18736), .n312(n312)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(82[5] 88[4])
    VLO i1 (.Z(GND_net));
    LUT4 i7459_2_lut_rep_433 (.A(count_beat[0]), .B(n4689), .Z(n18615)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i7459_2_lut_rep_433.init = 16'h8888;
    LUT4 i7991_2_lut_rep_622 (.A(count_note[1]), .B(count_note[2]), .Z(n18804)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i7991_2_lut_rep_622.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(count_note[1]), .B(count_note[2]), .C(count_note[4]), 
         .Z(n8_adj_1487)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i8172_3_lut_4_lut (.A(count_note[1]), .B(count_note[2]), .C(count_note[3]), 
         .D(count_note[4]), .Z(n13027)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i8172_3_lut_4_lut.init = 16'hf800;
    LUT4 i8009_2_lut_3_lut_3_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n22_adj_1459)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i8009_2_lut_3_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut_adj_62 (.A(count_note[1]), .B(count_note[2]), .C(count_note[4]), 
         .Z(n4)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i1_2_lut_3_lut_adj_62.init = 16'hf7f7;
    FD1S3AX count_beat_i4_2224__i1 (.D(n29_adj_1480), .CK(clk__inv), .Q(count_beat[1]));   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam count_beat_i4_2224__i1.GSR = "DISABLED";
    LUT4 i7998_2_lut_3_lut_3_lut_3_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n22_adj_1442)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i7998_2_lut_3_lut_3_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i8164_2_lut_3_lut_3_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[0]), .D(count_note[3]), .Z(n14_adj_1460)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i8164_2_lut_3_lut_3_lut_4_lut.init = 16'hff7f;
    FD1S3AX count_beat_i4_2224__i2 (.D(n28), .CK(clk__inv), .Q(count_beat[2]));   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam count_beat_i4_2224__i2.GSR = "DISABLED";
    FD1S3AX count_beat_i4_2224__i3 (.D(n27), .CK(clk__inv), .Q(count_beat[3]));   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam count_beat_i4_2224__i3.GSR = "DISABLED";
    FD1S3AX count_beat_i4_2224__i4 (.D(n26_adj_1479), .CK(clk__inv), .Q(count_beat[4]));   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam count_beat_i4_2224__i4.GSR = "DISABLED";
    FD1S3IX cnt_2220__i1 (.D(n132), .CK(clk__inv), .CD(n10969), .Q(cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_489_3_lut_4_lut (.A(count_note[1]), .B(count_note[2]), 
         .C(count_note[3]), .D(count_note[0]), .Z(n18671)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i1_2_lut_rep_489_3_lut_4_lut.init = 16'hf8f0;
    FD1S3IX cnt_2220__i2 (.D(n131), .CK(clk__inv), .CD(n10969), .Q(cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i2.GSR = "ENABLED";
    FD1S3IX cnt_2220__i3 (.D(n130), .CK(clk__inv), .CD(n10969), .Q(cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i3.GSR = "ENABLED";
    FD1S3IX cnt_2220__i4 (.D(n129), .CK(clk__inv), .CD(n10969), .Q(cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i4.GSR = "ENABLED";
    FD1S3IX cnt_2220__i5 (.D(n128), .CK(clk__inv), .CD(n10969), .Q(cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i5.GSR = "ENABLED";
    FD1S3IX cnt_2220__i6 (.D(n127), .CK(clk__inv), .CD(n10969), .Q(cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i6.GSR = "ENABLED";
    FD1S3IX cnt_2220__i7 (.D(n126), .CK(clk__inv), .CD(n10969), .Q(cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i7.GSR = "ENABLED";
    FD1S3IX cnt_2220__i8 (.D(n125), .CK(clk__inv), .CD(n10969), .Q(cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i8.GSR = "ENABLED";
    FD1S3IX cnt_2220__i9 (.D(n124), .CK(clk__inv), .CD(n10969), .Q(cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i9.GSR = "ENABLED";
    FD1S3IX cnt_2220__i10 (.D(n123), .CK(clk__inv), .CD(n10969), .Q(cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i10.GSR = "ENABLED";
    FD1S3IX cnt_2220__i11 (.D(n122), .CK(clk__inv), .CD(n10969), .Q(cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i11.GSR = "ENABLED";
    FD1S3IX cnt_2220__i12 (.D(n121), .CK(clk__inv), .CD(n10969), .Q(cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i12.GSR = "ENABLED";
    FD1S3IX cnt_2220__i13 (.D(n120), .CK(clk__inv), .CD(n10969), .Q(cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i13.GSR = "ENABLED";
    FD1S3IX cnt_2220__i14 (.D(n119), .CK(clk__inv), .CD(n10969), .Q(cnt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i14.GSR = "ENABLED";
    FD1S3IX cnt_2220__i15 (.D(n118), .CK(clk__inv), .CD(n10969), .Q(cnt[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i15.GSR = "ENABLED";
    FD1S3IX cnt_2220__i16 (.D(n117), .CK(clk__inv), .CD(n10969), .Q(cnt[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i16.GSR = "ENABLED";
    FD1S3IX cnt_2220__i17 (.D(n116), .CK(clk__inv), .CD(n10969), .Q(cnt[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i17.GSR = "ENABLED";
    FD1S3IX cnt_2220__i18 (.D(n115_adj_1502), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i18.GSR = "ENABLED";
    FD1S3IX cnt_2220__i19 (.D(n114_adj_1501), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i19.GSR = "ENABLED";
    FD1S3IX cnt_2220__i20 (.D(n113_adj_1500), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i20.GSR = "ENABLED";
    FD1S3IX cnt_2220__i21 (.D(n112_adj_1499), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i21.GSR = "ENABLED";
    FD1S3IX cnt_2220__i22 (.D(n111_adj_1498), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i22.GSR = "ENABLED";
    FD1S3IX cnt_2220__i23 (.D(n110_adj_1497), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i23.GSR = "ENABLED";
    FD1S3IX cnt_2220__i24 (.D(n109_adj_1496), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i24.GSR = "ENABLED";
    FD1S3IX cnt_2220__i25 (.D(n108_adj_1495), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i25.GSR = "ENABLED";
    FD1S3IX cnt_2220__i26 (.D(n107_adj_1494), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i26.GSR = "ENABLED";
    FD1S3IX cnt_2220__i27 (.D(n106_adj_1493), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i27.GSR = "ENABLED";
    FD1S3IX cnt_2220__i28 (.D(n105_adj_1492), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i28.GSR = "ENABLED";
    FD1S3IX cnt_2220__i29 (.D(n104_adj_1491), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[29])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i29.GSR = "ENABLED";
    FD1S3IX cnt_2220__i30 (.D(n103_adj_1490), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[30])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i30.GSR = "ENABLED";
    FD1S3IX cnt_2220__i31 (.D(n102_adj_1489), .CK(clk__inv), .CD(n10969), 
            .Q(cnt[31])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220__i31.GSR = "ENABLED";
    PFUMX mux_617_Mux_0_i109 (.BLUT(n101_adj_1511), .ALUT(n108_adj_1510), 
          .C0(count_note[4]), .Z(n109_adj_1509));
    L6MUX21 i11829 (.D0(n17190), .D1(n17197), .SD(count_note[6]), .Z(n17120));
    L6MUX21 i11826 (.D0(n17181), .D1(n17184), .SD(count_note[6]), .Z(n17117));
    L6MUX21 i11841 (.D0(n17130), .D1(n17131), .SD(count_note[6]), .Z(n17132));
    LUT4 i7943_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n86), 
         .Z(n106)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7943_2_lut_3_lut.init = 16'hd0d0;
    L6MUX21 i11927 (.D0(n17155), .D1(n17158), .SD(count_note[6]), .Z(n17218));
    key_U14 u_key_8 (.clk_N_168(clk_N_168), .\key_flag[7] (key_flag[7]), 
            .key_c_7(key_c_7), .\key_value[7] (key_value[7]), .GND_net(GND_net), 
            .n18756(n18756), .n18770(n18770), .n18758(n18758), .n37(n37), 
            .n34(n34), .\cycle_17__N_740[10] (cycle_17__N_740[10]), .n19846(n19846), 
            .\cycle_17__N_663[10] (cycle_17__N_663[10]), .n18815(n18815), 
            .\key_flag[8] (key_flag[8]), .\key_value[8] (key_value[8]), 
            .n18685(n18685), .\key_flag[6] (key_flag[6]), .\key_value[6] (key_value[6]), 
            .n18708(n18708), .n456(n456), .n3800(n3800), .n464(n464), 
            .n3815(n3815)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(107[5] 113[4])
    PFUMX i21 (.BLUT(n6_adj_1488), .ALUT(n8_adj_1487), .C0(count_note[6]), 
          .Z(n10));
    L6MUX21 i11839 (.D0(n17126), .D1(n17127), .SD(count_note[5]), .Z(n17130));
    L6MUX21 i11840 (.D0(n17128), .D1(n17129), .SD(count_note[5]), .Z(n17131));
    L6MUX21 i11847 (.D0(n17136), .D1(n17137), .SD(count_note[5]), .Z(n17138));
    L6MUX21 i11854 (.D0(n17143), .D1(n17144), .SD(count_note[5]), .Z(n17145));
    L6MUX21 i11857 (.D0(n17146), .D1(n17147), .SD(count_note[5]), .Z(n17148));
    L6MUX21 i11864 (.D0(n17153), .D1(n17154), .SD(count_note[5]), .Z(n17155));
    L6MUX21 i11867 (.D0(n17156), .D1(n17157), .SD(count_note[5]), .Z(n17158));
    L6MUX21 i11873 (.D0(n17162), .D1(n17163), .SD(count_note[5]), .Z(n17164));
    key_U27 u_key_10 (.GND_net(GND_net), .clk_N_168(clk_N_168), .\key_flag[9] (key_flag[9]), 
            .key_c_9(key_c_9), .\key_value[9] (key_value[9]), .n18768(n18768), 
            .\key_flag[8] (key_flag[8]), .\key_value[8] (key_value[8]), 
            .n9654(n9654), .\rom2[0] (rom2[0]), .n18771(n18771), .n17235(n17235), 
            .n6(n6_adj_1446), .n5(n5_adj_1445), .n911(n911)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(124[5] 130[4])
    L6MUX21 i11880 (.D0(n17169), .D1(n17170), .SD(count_note[5]), .Z(n17171));
    L6MUX21 i11890 (.D0(n17179), .D1(n17180), .SD(count_note[5]), .Z(n17181));
    L6MUX21 i11893 (.D0(n17182), .D1(n17183), .SD(count_note[5]), .Z(n17184));
    L6MUX21 i11896 (.D0(n17185), .D1(n17186), .SD(count_note[5]), .Z(n17187));
    L6MUX21 i11899 (.D0(n17188), .D1(n17189), .SD(count_note[5]), .Z(n17190));
    key_U26 u_key_11 (.clk_N_168(clk_N_168), .\key_flag[10] (key_flag[10]), 
            .key_c_10(key_c_10), .\key_value[10] (key_value[10]), .GND_net(GND_net), 
            .n18771(n18771), .n18761(n18761), .n344(n344), .n18763(n18763), 
            .n407(n407), .n9654(n9654), .n312(n312), .n18709(n18709), 
            .n417(n417), .n18768(n18768), .n321(n321), .n405(n405), 
            .\key_flag[11] (key_flag[11]), .\key_value[11] (key_value[11]), 
            .n16909(n16909), .n6(n6_adj_1446), .n18813(n18813), .n18719(n18719), 
            .\key_value[9] (key_value[9]), .\key_flag[9] (key_flag[9]), 
            .n18667(n18667)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(132[5] 138[4])
    L6MUX21 i11906 (.D0(n17195), .D1(n17196), .SD(count_note[5]), .Z(n17197));
    L6MUX21 i11913 (.D0(n17202), .D1(n17203), .SD(count_note[5]), .Z(n17204));
    L6MUX21 i11916 (.D0(n17205), .D1(n17206), .SD(count_note[5]), .Z(n17207));
    L6MUX21 i11926 (.D0(n17215), .D1(n17216), .SD(count_note[5]), .Z(n17217));
    key_U25 u_key_12 (.clk_N_168(clk_N_168), .\key_flag[11] (key_flag[11]), 
            .key_c_11(key_c_11), .\key_value[11] (key_value[11]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(140[5] 146[4])
    L6MUX21 i11936 (.D0(n17225), .D1(n17226), .SD(count_note[5]), .Z(n17227));
    key_U20 u_key_2 (.clk_N_168(clk_N_168), .\key_flag[1] (key_flag[1]), 
            .key_c_1(key_c_1), .\key_value[1] (key_value[1]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(57[5] 63[4])
    PFUMX i11897 (.BLUT(n7_adj_1503), .ALUT(n14_adj_1460), .C0(count_note[4]), 
          .Z(n17188));
    PFUMX i11894 (.BLUT(n70_adj_1505), .ALUT(n77_adj_1504), .C0(count_note[4]), 
          .Z(n17185));
    PFUMX i11891 (.BLUT(n38_adj_1462), .ALUT(n10407), .C0(count_note[4]), 
          .Z(n17182));
    key_U24 u_key_13 (.clk_N_168(clk_N_168), .\key_flag[12] (key_flag[12]), 
            .key_c_12(key_c_12), .\key_value[12] (key_value[12]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(148[5] 154[4])
    PFUMX i11871 (.BLUT(n13008), .ALUT(n14_adj_1466), .C0(count_note[4]), 
          .Z(n17162));
    LUT4 mux_674_Mux_2_i109_then_4_lut (.A(count_note[4]), .B(count_note[3]), 
         .C(count_note[1]), .D(count_note[2]), .Z(n18840)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C)+!B ((D)+!C)))) */ ;
    defparam mux_674_Mux_2_i109_then_4_lut.init = 16'h0416;
    PFUMX i11845 (.BLUT(n7_adj_1441), .ALUT(n14), .C0(count_note[4]), 
          .Z(n17136));
    LUT4 i7944_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n85), 
         .Z(n105)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7944_2_lut_3_lut.init = 16'hd0d0;
    key_U13 u_key_9 (.clk_N_168(clk_N_168), .\key_flag[8] (key_flag[8]), 
            .key_c_8(key_c_8), .\key_value[8] (key_value[8]), .GND_net(GND_net), 
            .n18755(n18755), .\rom2[0] (rom2[0]), .n18815(n18815), .n17234(n17234), 
            .n18770(n18770), .n5(n5), .n464(n464), .n6(n6_adj_1446), 
            .n5_adj_2(n5_adj_1447), .n907(n907), .n18768(n18768), .n16917(n16917)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(116[5] 122[4])
    LUT4 i7997_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n22_adj_1463)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i7997_4_lut_4_lut_4_lut.init = 16'h70c0;
    LUT4 mux_674_Mux_2_i109_else_4_lut (.A(count_note[4]), .B(count_note[3]), 
         .C(count_note[1]), .D(count_note[2]), .Z(n18839)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam mux_674_Mux_2_i109_else_4_lut.init = 16'h4324;
    PFUMX i11835 (.BLUT(n7_adj_1486), .ALUT(n14_adj_1485), .C0(count_note[4]), 
          .Z(n17126));
    LUT4 i15_2_lut_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), .C(count_note[3]), 
         .D(count_note[2]), .Z(n16773)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i15_2_lut_3_lut_4_lut.init = 16'hf087;
    key_U21 u_key_1 (.GND_net(GND_net), .\key_value[0] (key_value[0]), .clk_N_168(clk_N_168), 
            .key_c_0(key_c_0), .\key_flag[0] (key_flag[0]), .n5(n5), .n18721(n18721), 
            .n18724(n18724), .n9292(n9292), .n18644(n18644), .n6(n6), 
            .n5_adj_1(n5_adj_1447), .n18713(n18713), .n19846(n19846), 
            .n18680(n18680), .n18679(n18679), .n18722(n18722), .n18725(n18725), 
            .n18649(n18649), .n18652(n18652)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(48[5] 54[4])
    LUT4 mux_617_Mux_4_i14_4_lut_4_lut_3_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n14_adj_1485)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_4_i14_4_lut_4_lut_3_lut_4_lut.init = 16'h0778;
    LUT4 mux_674_Mux_1_i109_then_4_lut (.A(count_note[4]), .B(count_note[3]), 
         .C(count_note[1]), .D(count_note[2]), .Z(n18843)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A !((C+(D))+!B))) */ ;
    defparam mux_674_Mux_1_i109_then_4_lut.init = 16'h5771;
    LUT4 i2_3_lut_4_lut_4_lut (.A(count_note[0]), .B(n18804), .C(n16847), 
         .D(count_note[3]), .Z(n16854)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 mux_674_Mux_1_i109_else_4_lut (.A(count_note[4]), .B(count_note[3]), 
         .C(count_note[1]), .D(count_note[2]), .Z(n18842)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C (D))+!B !(C+!(D))))) */ ;
    defparam mux_674_Mux_1_i109_else_4_lut.init = 16'h1457;
    LUT4 i10423_2_lut_3_lut_4_lut_4_lut (.A(count_beat[0]), .B(n4689), .C(n18760), 
         .D(count_beat[1]), .Z(n29_adj_1480)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A !(B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i10423_2_lut_3_lut_4_lut_4_lut.init = 16'h4c80;
    LUT4 i39_then_4_lut (.A(count_note[4]), .B(count_note[3]), .C(count_note[1]), 
         .D(count_note[2]), .Z(n18846)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B ((D)+!C)+!B !(C (D))))) */ ;
    defparam i39_then_4_lut.init = 16'h4737;
    LUT4 i39_else_4_lut (.A(count_note[4]), .B(count_note[3]), .C(count_note[1]), 
         .D(count_note[2]), .Z(n18845)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B (D)+!B (C (D))))) */ ;
    defparam i39_else_4_lut.init = 16'h2357;
    LUT4 i5892_3_lut_rep_630 (.A(count_note[0]), .B(count_note[1]), .C(count_note[2]), 
         .D(count_note[3]), .Z(n18812)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i5892_3_lut_rep_630.init = 16'hff80;
    LUT4 i8189_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n108_adj_1510)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i8189_3_lut_4_lut_4_lut.init = 16'h0013;
    LUT4 i11923_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17214)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B ((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11923_3_lut_4_lut_4_lut_4_lut.init = 16'h8630;
    LUT4 i11921_3_lut_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17212)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A (B (C+(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11921_3_lut_3_lut_4_lut_4_lut.init = 16'h1186;
    LUT4 mux_617_Mux_3_i60_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n60_adj_1507)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_3_i60_3_lut_4_lut_4_lut.init = 16'h79cf;
    LUT4 i11900_3_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n17191)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A (B (C+(D))+!B !(C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11900_3_lut_4_lut_4_lut.init = 16'hcf79;
    LUT4 mux_617_Mux_2_i29_3_lut_4_lut_4_lut_4_lut (.A(count_note[0]), .B(count_note[1]), 
         .C(count_note[2]), .D(count_note[3]), .Z(n29_adj_1465)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_2_i29_3_lut_4_lut_4_lut_4_lut.init = 16'haf83;
    TSALL TSALL_INST (.TSALL(GND_net));
    PFUMX i11836 (.BLUT(n22_adj_1484), .ALUT(n13024), .C0(count_note[4]), 
          .Z(n17127));
    PFUMX i11837 (.BLUT(n38_adj_1483), .ALUT(n45_adj_1482), .C0(count_note[4]), 
          .Z(n17128));
    LUT4 i7945_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n84), 
         .Z(n104)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7945_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i11834_3_lut (.A(n17123), .B(n17124), .C(count_note[7]), .Z(beat_4__N_40[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11834_3_lut.init = 16'hcaca;
    LUT4 i11833_3_lut (.A(n17227), .B(n18841), .C(count_note[6]), .Z(n17124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11833_3_lut.init = 16'hcaca;
    LUT4 i11831_3_lut (.A(n17120), .B(n17121), .C(count_note[7]), .Z(beat_4__N_40[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11831_3_lut.init = 16'hcaca;
    key_U15 u_key_7 (.clk_N_168(clk_N_168), .\key_flag[6] (key_flag[6]), 
            .key_c_6(key_c_6), .\key_value[6] (key_value[6]), .GND_net(GND_net), 
            .n18720(n18720), .n18754(n18754), .n18815(n18815), .n18654(n18654), 
            .n18735(n18735), .n18655(n18655), .n6(n6_adj_1443), .n18813(n18813), 
            .n18677(n18677), .n18747(n18747), .n12156(n12156), .n456(n456), 
            .\rom2[1] (rom2[1]), .n18597(n18597), .n18755(n18755), .n18668(n18668)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(98[5] 104[4])
    LUT4 i11830_3_lut (.A(n17204), .B(n18844), .C(count_note[6]), .Z(n17121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11830_3_lut.init = 16'hcaca;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 n18443_bdd_3_lut_12700 (.A(n18443), .B(n18837), .C(count_note[3]), 
         .Z(n18444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n18443_bdd_3_lut_12700.init = 16'hcaca;
    PFUMX i11846 (.BLUT(n22_adj_1444), .ALUT(n10403), .C0(count_note[4]), 
          .Z(n17137));
    LUT4 i7936_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n93), 
         .Z(n113)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7936_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_617_Mux_4_i127_4_lut (.A(n17132), .B(n94), .C(count_note[7]), 
         .D(count_note[6]), .Z(note_5__N_45[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_4_i127_4_lut.init = 16'h0aca;
    LUT4 mux_617_Mux_4_i94_4_lut (.A(n17230), .B(n92_adj_1474), .C(count_note[5]), 
         .D(count_note[4]), .Z(n94)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_4_i94_4_lut.init = 16'hca0a;
    LUT4 i7935_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n94_adj_1477), 
         .Z(n114)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7935_2_lut_3_lut.init = 16'hd0d0;
    PFUMX i11852 (.BLUT(n17139), .ALUT(n17140), .C0(count_note[4]), .Z(n17143));
    LUT4 i11828_3_lut (.A(n17117), .B(n17118), .C(count_note[7]), .Z(note_5__N_45[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11828_3_lut.init = 16'hcaca;
    LUT4 i11827_4_lut (.A(n17187), .B(n18774), .C(count_note[6]), .D(n4), 
         .Z(n17118)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i11827_4_lut.init = 16'hfaca;
    key_U16 u_key_6 (.clk_N_168(clk_N_168), .\key_flag[5] (key_flag[5]), 
            .key_c_5(key_c_5), .\key_value[5] (key_value[5]), .GND_net(GND_net), 
            .n18754(n18754), .\key_value[4] (key_value[4]), .\key_flag[4] (key_flag[4]), 
            .n18706(n18706), .n6(n6_adj_1443), .n5(n5_adj_1445), .n895(n895)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(90[5] 96[4])
    LUT4 i11960_3_lut (.A(n17249), .B(n17250), .C(count_note[7]), .Z(note_5__N_45[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11960_3_lut.init = 16'hcaca;
    PFUMX i11853 (.BLUT(n17141), .ALUT(n17142), .C0(count_note[4]), .Z(n17144));
    LUT4 i11959_3_lut (.A(n18462), .B(n18847), .C(count_note[6]), .Z(n17250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11959_3_lut.init = 16'hcaca;
    LUT4 i10430_2_lut_3_lut_4_lut (.A(n18760), .B(n18615), .C(n8_adj_1478), 
         .D(n18614), .Z(n28)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i10430_2_lut_3_lut_4_lut.init = 16'h78f0;
    PFUMX i11855 (.BLUT(n70), .ALUT(n77), .C0(count_note[4]), .Z(n17146));
    FD1P3AX stat_71_rep_637 (.D(n17430), .SP(VCC_net), .CK(clk_N_168), 
            .Q(n19846)) /* synthesis lse_init_val=0 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(196[7] 205[5])
    defparam stat_71_rep_637.GSR = "ENABLED";
    LUT4 i11929_3_lut (.A(n17218), .B(n17219), .C(count_note[7]), .Z(note_5__N_45[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11929_3_lut.init = 16'hcaca;
    LUT4 i11928_4_lut (.A(n18444), .B(count_note[3]), .C(count_note[6]), 
         .D(n16_adj_1439), .Z(n17219)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam i11928_4_lut.init = 16'h3a0a;
    PFUMX i11856 (.BLUT(n10405), .ALUT(n92_adj_1512), .C0(count_note[4]), 
          .Z(n17147));
    PFUMX i11862 (.BLUT(n17149), .ALUT(n17150), .C0(count_note[4]), .Z(n17153));
    PFUMX i11863 (.BLUT(n17151), .ALUT(n17152), .C0(count_note[4]), .Z(n17154));
    CCU2D cnt_2220_add_4_33 (.A0(cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15798), .S0(n102_adj_1489));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_33.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_33.INIT1 = 16'h0000;
    defparam cnt_2220_add_4_33.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_33.INJECT1_1 = "NO";
    LUT4 LessThan_51_i7_2_lut_rep_544 (.A(count_beat[3]), .B(beat[3]), .Z(n18726)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(242[8:25])
    defparam LessThan_51_i7_2_lut_rep_544.init = 16'h6666;
    LUT4 LessThan_51_i6_3_lut_3_lut (.A(count_beat[3]), .B(beat[3]), .C(beat[2]), 
         .Z(n6_adj_1451)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(242[8:25])
    defparam LessThan_51_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 LessThan_51_i9_2_lut_rep_545 (.A(count_beat[4]), .B(beat[4]), .Z(n18727)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(242[8:25])
    defparam LessThan_51_i9_2_lut_rep_545.init = 16'h6666;
    LUT4 i7939_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n90), 
         .Z(n110)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7939_2_lut_3_lut.init = 16'hd0d0;
    LUT4 LessThan_51_i8_3_lut_3_lut (.A(count_beat[4]), .B(beat[4]), .C(n6_adj_1451), 
         .Z(n8)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(242[8:25])
    defparam LessThan_51_i8_3_lut_3_lut.init = 16'hd4d4;
    PFUMX i11865 (.BLUT(n38_adj_1468), .ALUT(n45_adj_1469), .C0(count_note[4]), 
          .Z(n17156));
    PFUMX i11866 (.BLUT(n53), .ALUT(n60), .C0(count_note[4]), .Z(n17157));
    LUT4 i2_3_lut_4_lut (.A(count_note[2]), .B(count_note[3]), .C(count_note[5]), 
         .D(count_note[6]), .Z(n16859)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i2_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_548 (.A(count_note[5]), .B(count_note[6]), .Z(n18730)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i1_2_lut_rep_548.init = 16'h2222;
    PFUMX i11872 (.BLUT(n22_adj_1464), .ALUT(n29_adj_1465), .C0(count_note[4]), 
          .Z(n17163));
    LUT4 i1_2_lut_3_lut_4_lut_adj_63 (.A(count_note[5]), .B(count_note[6]), 
         .C(count_note[3]), .D(count_note[2]), .Z(n16869)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(518[2] 775[12])
    defparam i1_2_lut_3_lut_4_lut_adj_63.init = 16'h0002;
    FD1P3IX count_note_2222__i7 (.D(n38_adj_1457), .SP(clk_N_168_enable_533), 
            .CD(n10968), .CK(clk_N_168), .Q(count_note[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i7.GSR = "DISABLED";
    LUT4 i2_3_lut_3_lut (.A(count_note[0]), .B(count_note[7]), .C(n10), 
         .Z(beat_4__N_40[3])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i2_3_lut_3_lut.init = 16'h4040;
    PFUMX i11878 (.BLUT(n17165), .ALUT(n17166), .C0(count_note[4]), .Z(n17169));
    FD1P3IX count_note_2222__i6 (.D(n39), .SP(clk_N_168_enable_533), .CD(n10968), 
            .CK(clk_N_168), .Q(count_note[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i6.GSR = "DISABLED";
    PFUMX i11879 (.BLUT(n17167), .ALUT(n17168), .C0(count_note[4]), .Z(n17170));
    FD1P3IX count_note_2222__i5 (.D(n40_adj_1456), .SP(clk_N_168_enable_533), 
            .CD(n10968), .CK(clk_N_168), .Q(count_note[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i5.GSR = "DISABLED";
    LUT4 mux_617_Mux_1_i60_4_lut_4_lut (.A(count_note[2]), .B(count_note[3]), 
         .C(n18781), .D(n37_adj_1467), .Z(n60)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam mux_617_Mux_1_i60_4_lut_4_lut.init = 16'h7340;
    LUT4 i11882_4_lut_4_lut_4_lut (.A(count_note[2]), .B(count_note[0]), 
         .C(count_note[3]), .D(count_note[1]), .Z(n17173)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C+(D))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(256[5] 513[9])
    defparam i11882_4_lut_4_lut_4_lut.init = 16'ha0ad;
    FD1P3IX count_note_2222__i4 (.D(n41_adj_1455), .SP(clk_N_168_enable_533), 
            .CD(n10968), .CK(clk_N_168), .Q(count_note[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i4.GSR = "DISABLED";
    CCU2D cnt_2220_add_4_31 (.A0(cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15797), .COUT(n15798), .S0(n104_adj_1491), .S1(n103_adj_1490));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_31.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_31.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_31.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_31.INJECT1_1 = "NO";
    FD1P3AX beat_i0 (.D(beat_4__N_40[0]), .SP(clk_N_168_enable_534), .CK(clk_N_168), 
            .Q(beat[0]));   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam beat_i0.GSR = "DISABLED";
    FD1P3IX count_note_2222__i3 (.D(n42_adj_1454), .SP(clk_N_168_enable_533), 
            .CD(n10968), .CK(clk_N_168), .Q(count_note[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i3.GSR = "DISABLED";
    key_U19 u_key_3 (.clk_N_168(clk_N_168), .\key_flag[2] (key_flag[2]), 
            .key_c_2(key_c_2), .\key_value[2] (key_value[2]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(66[5] 72[4])
    PFUMX i11888 (.BLUT(n7_adj_1461), .ALUT(n16773), .C0(count_note[4]), 
          .Z(n17179));
    GSR GSR_INST (.GSR(rst_n_c));
    PFUMX i11889 (.BLUT(n22_adj_1463), .ALUT(n16860), .C0(count_note[4]), 
          .Z(n17180));
    PFUMX i11892 (.BLUT(n53_adj_1508), .ALUT(n60_adj_1507), .C0(count_note[4]), 
          .Z(n17183));
    PFUMX i11895 (.BLUT(n16896), .ALUT(n92), .C0(count_note[4]), .Z(n17186));
    LUT4 i7953_2_lut (.A(count_beat[2]), .B(n4689), .Z(n8_adj_1478)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(241[4] 251[7])
    defparam i7953_2_lut.init = 16'h8888;
    PFUMX i11898 (.BLUT(n22_adj_1459), .ALUT(n29_adj_1458), .C0(count_note[4]), 
          .Z(n17189));
    FD1P3IX count_note_2222__i2 (.D(n43), .SP(clk_N_168_enable_533), .CD(n10968), 
            .CK(clk_N_168), .Q(count_note[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i2.GSR = "DISABLED";
    FD1P3IX count_note_2222__i1 (.D(n44_adj_1453), .SP(clk_N_168_enable_533), 
            .CD(n10968), .CK(clk_N_168), .Q(count_note[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(247[24:39])
    defparam count_note_2222__i1.GSR = "DISABLED";
    LUT4 n16859_bdd_4_lut (.A(n16859), .B(n16869), .C(count_note[7]), 
         .D(count_note[1]), .Z(n18604)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n16859_bdd_4_lut.init = 16'hca00;
    PFUMX i11904 (.BLUT(n17191), .ALUT(n17192), .C0(count_note[4]), .Z(n17195));
    PFUMX i11905 (.BLUT(n17193), .ALUT(n17194), .C0(count_note[4]), .Z(n17196));
    CCU2D cnt_2220_add_4_29 (.A0(cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15796), .COUT(n15797), .S0(n106_adj_1493), .S1(n105_adj_1492));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_29.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_29.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_29.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_29.INJECT1_1 = "NO";
    FD1P3AX beat_i3 (.D(beat_4__N_40[3]), .SP(clk_N_168_enable_534), .CK(clk_N_168), 
            .Q(beat[3]));   // d:/fpga_project/lattice_diamond/piano/piano.v(517[7] 776[4])
    defparam beat_i3.GSR = "DISABLED";
    PFUMX i11911 (.BLUT(n17198), .ALUT(n17199), .C0(count_note[4]), .Z(n17202));
    CCU2D cnt_2220_add_4_27 (.A0(cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15795), .COUT(n15796), .S0(n108_adj_1495), .S1(n107_adj_1494));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_27.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_27.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_27.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_27.INJECT1_1 = "NO";
    key_U22 u_key_15 (.clk_N_168(clk_N_168), .\key_flag[14] (key_flag[14]), 
            .key_c_14(key_c_14), .\key_value[14] (key_value[14]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(164[5] 170[4])
    PFUMX i11912 (.BLUT(n17200), .ALUT(n17201), .C0(count_note[4]), .Z(n17203));
    CCU2D cnt_2220_add_4_25 (.A0(cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15794), .COUT(n15795), .S0(n110_adj_1497), .S1(n109_adj_1496));   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam cnt_2220_add_4_25.INIT0 = 16'hfaaa;
    defparam cnt_2220_add_4_25.INIT1 = 16'hfaaa;
    defparam cnt_2220_add_4_25.INJECT1_0 = "NO";
    defparam cnt_2220_add_4_25.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_64 (.A(n19846), .B(rom2[3]), .C(n17135), .D(n58), 
         .Z(en_1__N_194)) /* synthesis lut_function=(A+!(B ((D)+!C)+!B !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(196[7] 205[5])
    defparam i1_4_lut_adj_64.init = 16'hbafa;
    LUT4 i12350_2_lut (.A(cnt[0]), .B(n10216), .Z(n10969)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(228[12:17])
    defparam i12350_2_lut.init = 16'h2222;
    PFUMX i11914 (.BLUT(n7), .ALUT(n14_adj_1440), .C0(count_note[4]), 
          .Z(n17205));
    key_U18 u_key_4 (.clk_N_168(clk_N_168), .\key_flag[3] (key_flag[3]), 
            .key_c_3(key_c_3), .\key_value[3] (key_value[3]), .GND_net(GND_net), 
            .n18736(n18736), .n6(n6_adj_1443), .n18814(n18814), .n887(n887), 
            .\rom2[1] (rom2[1]), .n18754(n18754), .n18598(n18598), .\key_flag[2] (key_flag[2]), 
            .\key_value[2] (key_value[2]), .n18707(n18707), .n18747(n18747), 
            .n18758(n18758), .n444(n444), .\key_value[4] (key_value[4]), 
            .\key_flag[4] (key_flag[4]), .n18696(n18696)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(74[5] 80[4])
    clk_pll u_clk_pll (.sys_clk_c(sys_clk_c), .clk(clk), .GND_net(GND_net), 
            .clk_N_168(clk_N_168)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(31[9] 34[5])
    PFUMX i11915 (.BLUT(n22_adj_1442), .ALUT(n29), .C0(count_note[4]), 
          .Z(n17206));
    PFUMX i11924 (.BLUT(n17211), .ALUT(n17212), .C0(count_note[4]), .Z(n17215));
    LUT4 i12347_3_lut (.A(n19846), .B(clk_beat), .C(n201), .Z(clk_N_168_enable_533)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(240[3] 252[9])
    defparam i12347_3_lut.init = 16'h0808;
    LUT4 i12356_4_lut (.A(clk_N_168_enable_533), .B(n13027), .C(n16847), 
         .D(count_note[5]), .Z(n10968)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i12356_4_lut.init = 16'ha080;
    PFUMX i11925 (.BLUT(n17213), .ALUT(n17214), .C0(count_note[4]), .Z(n17216));
    PFUMX i11934 (.BLUT(n17221), .ALUT(n17222), .C0(count_note[4]), .Z(n17225));
    PFUMX i11935 (.BLUT(n17223), .ALUT(n17224), .C0(count_note[4]), .Z(n17226));
    LUT4 i4_4_lut (.A(n7_adj_1448), .B(n18730), .C(count_note[7]), .D(count_note[4]), 
         .Z(beat_4__N_40[0])) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0800;
    PFUMX LessThan_51_i10 (.BLUT(n4_adj_1452), .ALUT(n8), .C0(n17020), 
          .Z(n201));
    PFUMX i11939 (.BLUT(n17228), .ALUT(n17229), .C0(count_note[4]), .Z(n17230));
    LUT4 i7942_2_lut_3_lut (.A(n3759), .B(CNT_17__N_703[18]), .C(n87), 
         .Z(n107)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i7942_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i12365_4_lut (.A(n18727), .B(n18726), .C(count_beat[2]), .D(beat[2]), 
         .Z(n17020)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(242[8:25])
    defparam i12365_4_lut.init = 16'heffe;
    key_U23 u_key_14 (.clk_N_168(clk_N_168), .\key_flag[13] (key_flag[13]), 
            .key_c_13(key_c_13), .\key_value[13] (key_value[13]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(156[5] 162[4])
    LUT4 i12269_2_lut (.A(cnt[0]), .B(n10216), .Z(clk_beat_N_126)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(233[5:17])
    defparam i12269_2_lut.init = 16'h1111;
    PFUMX i11838 (.BLUT(n16868), .ALUT(n16865), .C0(count_note[4]), .Z(n17129));
    
endmodule
//
// Verilog Description of module speaker
//

module speaker (GND_net, \PWM_in_12__N_452[2] , \PWM_in_12__N_452[3] , 
            \data_out1[0] , \data_out2[0] , \PWM_in_12__N_452[1] , n9292, 
            \rom1_4__N_338[0] , \rom2[0] , clk_N_168, n19846, \key_value[4] , 
            n28, stat, \yinjie_box_2__N_394[0] , \yinjie_box_2__N_394[1] , 
            \key_value[10] , n18598, n18597, n18644, \rom2[1] , \rom2[3] , 
            \key_value[5] , \key_value[1] , \key_value[12] , \key_value[11] , 
            \key_flag[8] , \key_flag[0] , n5, n18808, \note[0] , \note[1] , 
            n18737, n7, n18807, n18803, n18307, n6, n18610, \cycle_17__N_663[17] , 
            n18719, n911, n907, n895, n18677, n887, n891, n18713, 
            n456, n444, n11464, n18676, n436, n18679, n5_adj_11, 
            \key_flag[9] , \key_flag[10] , \note[4] , \note[3] , \note[2] , 
            n18747, n18754, \key_flag[1] , \key_flag[2] , n18722, 
            n12156, n18724, n18720, n18813, n6_adj_12, n18763, n18761, 
            n16917, n9654, n16909, n10160, n406, n18755, n18667, 
            n410, n18815, n31, n321, n6_adj_13, pwm_out2_c, \cycle_17__N_663[7] , 
            n14_adj_14, n3, \cycle_17__N_740[12] , n18772, n3_adj_15, 
            \cycle_17__N_740[11] , n7_adj_16, n18734, \key_value[7] , 
            \key_value[9] , n18758, \key_value[8] , \key_flag[11] , 
            n18771, n18814, n18768, n18620, n5_adj_17, \key_flag[12] , 
            n18709, n18770, \key_value[0] , n18685, n18619, n16876, 
            clk_N_168_enable_512, n18736, n18735, n18725, n247, n18708, 
            n9, n331, n415, n18651, n18308, n18850, \key_value[2] , 
            \key_value[3] , \key_value[6] , n26_adj_18, \cycle_17__N_663[2] , 
            n10337, n18707, n269, n22_adj_19, n18769, n16920, n18612, 
            n16959, n18623, n417, \cycle_17__N_740[1] , n18697, \cycle_17__N_740[14] , 
            n19_adj_20, n17110, n12983, n9757, n17135, \PWM_in_12__N_452[12] , 
            n37, n464, \key_flag[3] , \key_flag[5] , \key_flag[6] , 
            n18756, n34, en_1__N_194, n18606, n18721, n18668, n3815, 
            n3830, n3800, \key_flag[4] , \key_flag[7] , n18684, n18682, 
            n16828, n18706, n16888, n18616, \cycle_17__N_740[3] , 
            n414, \cycle_17__N_740[4] , \cycle_17__N_740[16] , n405, 
            \cycle_17__N_740[13] , n262, \cycle_17__N_740[9] , \PWM_in_12__N_452[10] , 
            \PWM_in_12__N_452[11] , \PWM_in_12__N_452[8] , \PWM_in_12__N_452[9] , 
            \PWM_in_12__N_452[6] , \PWM_in_12__N_452[7] , \PWM_in_12__N_452[4] , 
            \PWM_in_12__N_452[5] , n58, n351, n18655, n18680, clk_N_168_enable_507, 
            clk_N_168_enable_518, n17234, n17235, n18785, n18784, 
            n18757, n18717, n19839, \fcw_r_15__N_495[11] , \fcw_r_15__N_495[5] , 
            n8147, n8146, yinjie, clk__inv, \fcw_r_15__N_495[9] , 
            clk, rst_n_c, key_pa_c, \fcw_r_15__N_495[10] , \fcw_r_15__N_495[6] , 
            \fcw_r_15__N_495[8] , n18690, n10972, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \PWM_in_12__N_452[2] ;
    output \PWM_in_12__N_452[3] ;
    output \data_out1[0] ;
    output \data_out2[0] ;
    output \PWM_in_12__N_452[1] ;
    input n9292;
    input \rom1_4__N_338[0] ;
    output \rom2[0] ;
    input clk_N_168;
    input n19846;
    input \key_value[4] ;
    input [12:0]n28;
    input stat;
    output \yinjie_box_2__N_394[0] ;
    output \yinjie_box_2__N_394[1] ;
    input \key_value[10] ;
    input n18598;
    input n18597;
    input n18644;
    output \rom2[1] ;
    output \rom2[3] ;
    input \key_value[5] ;
    input \key_value[1] ;
    input \key_value[12] ;
    input \key_value[11] ;
    input \key_flag[8] ;
    input \key_flag[0] ;
    output n5;
    output n18808;
    input \note[0] ;
    input \note[1] ;
    output n18737;
    output n7;
    output n18807;
    input n18803;
    output n18307;
    output n6;
    output n18610;
    output \cycle_17__N_663[17] ;
    input n18719;
    input n911;
    input n907;
    input n895;
    input n18677;
    input n887;
    input n891;
    input n18713;
    input n456;
    input n444;
    input n11464;
    output n18676;
    output n436;
    input n18679;
    output n5_adj_11;
    input \key_flag[9] ;
    input \key_flag[10] ;
    input \note[4] ;
    input \note[3] ;
    input \note[2] ;
    output n18747;
    input n18754;
    input \key_flag[1] ;
    input \key_flag[2] ;
    output n18722;
    output n12156;
    output n18724;
    input n18720;
    output n18813;
    output n6_adj_12;
    output n18763;
    output n18761;
    input n16917;
    input n9654;
    input n16909;
    output n10160;
    output n406;
    input n18755;
    input n18667;
    output n410;
    input n18815;
    input n31;
    output n321;
    output n6_adj_13;
    output pwm_out2_c;
    output \cycle_17__N_663[7] ;
    input n14_adj_14;
    output n3;
    output \cycle_17__N_740[12] ;
    input n18772;
    output n3_adj_15;
    output \cycle_17__N_740[11] ;
    output n7_adj_16;
    input n18734;
    input \key_value[7] ;
    input \key_value[9] ;
    output n18758;
    input \key_value[8] ;
    input \key_flag[11] ;
    input n18771;
    output n18814;
    input n18768;
    output n18620;
    output n5_adj_17;
    input \key_flag[12] ;
    output n18709;
    output n18770;
    input \key_value[0] ;
    input n18685;
    input n18619;
    input n16876;
    output clk_N_168_enable_512;
    input n18736;
    input n18735;
    output n18725;
    output n247;
    input n18708;
    output n9;
    input n331;
    output n415;
    input n18651;
    output n18308;
    input n18850;
    input \key_value[2] ;
    input \key_value[3] ;
    input \key_value[6] ;
    input n26_adj_18;
    output \cycle_17__N_663[2] ;
    output n10337;
    input n18707;
    output n269;
    output n22_adj_19;
    input n18769;
    output n16920;
    output n18612;
    output n16959;
    output n18623;
    input n417;
    output \cycle_17__N_740[1] ;
    output n18697;
    output \cycle_17__N_740[14] ;
    output n19_adj_20;
    output n17110;
    output n12983;
    output n9757;
    output n17135;
    output \PWM_in_12__N_452[12] ;
    input n37;
    input n464;
    input \key_flag[3] ;
    input \key_flag[5] ;
    input \key_flag[6] ;
    input n18756;
    output n34;
    input en_1__N_194;
    output n18606;
    input n18721;
    input n18668;
    input n3815;
    output n3830;
    output n3800;
    input \key_flag[4] ;
    input \key_flag[7] ;
    output n18684;
    output n18682;
    input n16828;
    input n18706;
    input n16888;
    output n18616;
    output \cycle_17__N_740[3] ;
    input n414;
    output \cycle_17__N_740[4] ;
    output \cycle_17__N_740[16] ;
    input n405;
    output \cycle_17__N_740[13] ;
    input n262;
    output \cycle_17__N_740[9] ;
    output \PWM_in_12__N_452[10] ;
    output \PWM_in_12__N_452[11] ;
    output \PWM_in_12__N_452[8] ;
    output \PWM_in_12__N_452[9] ;
    output \PWM_in_12__N_452[6] ;
    output \PWM_in_12__N_452[7] ;
    output \PWM_in_12__N_452[4] ;
    output \PWM_in_12__N_452[5] ;
    output n58;
    output n351;
    input n18655;
    input n18680;
    output clk_N_168_enable_507;
    output clk_N_168_enable_518;
    input n17234;
    input n17235;
    output n18785;
    output n18784;
    input n18757;
    input n18717;
    input n19839;
    input \fcw_r_15__N_495[11] ;
    input \fcw_r_15__N_495[5] ;
    input n8147;
    input n8146;
    input [2:0]yinjie;
    output clk__inv;
    input \fcw_r_15__N_495[9] ;
    input clk;
    input rst_n_c;
    input key_pa_c;
    input \fcw_r_15__N_495[10] ;
    input \fcw_r_15__N_495[6] ;
    input \fcw_r_15__N_495[8] ;
    input n18690;
    input n10972;
    input VCC_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire clk /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    
    wire n15477;
    wire [11:0]data_out1;   // d:/fpga_project/lattice_diamond/piano/speaker.v(21[14:23])
    wire [11:0]data_out2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(22[17:26])
    
    wire n15478;
    wire [4:0]rom1;   // d:/fpga_project/lattice_diamond/piano/speaker.v(18[12:16])
    
    wire rom1_4__N_289, rom2_4__N_297;
    wire [4:0]rom2_4__N_397;
    wire [24:0]u_count1;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [24:0]u_count1_24__N_142;
    wire [24:0]count_24__N_543;
    wire [24:0]n52;
    wire [13:0]PWM_DDS_accumulator;   // d:/fpga_project/lattice_diamond/piano/speaker.v(23[16:35])
    
    wire pwm_out2_N_125;
    wire [12:0]n4943;
    wire [12:0]PWM_in;   // d:/fpga_project/lattice_diamond/piano/speaker.v(20[13:19])
    wire [18:0]fcw_r_15__N_527;
    wire [2:0]yinjie_box;   // d:/fpga_project/lattice_diamond/piano/speaker.v(24[12:22])
    wire [24:0]count_24__N_543_adj_1400;
    wire [24:0]n52_adj_1401;
    
    wire n18851, n18852, n3086, n18599;
    wire [3:0]n3836;
    
    wire n18622, n16818, n16916, n15957, n18643, n16903;
    wire [4:0]rom2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(18[27:31])
    
    wire n18621, n16823, n16930, n15938;
    wire [24:0]count_24__N_543_adj_1402;
    wire [24:0]n52_adj_1403;
    wire [24:0]count_24__N_543_adj_1404;
    wire [24:0]n52_adj_1405;
    wire [24:0]count1;   // d:/fpga_project/lattice_diamond/piano/speaker.v(11[15:21])
    wire [24:0]count3;   // d:/fpga_project/lattice_diamond/piano/speaker.v(11[53:59])
    wire [24:0]n3371;
    
    wire n18592, n18591, n17004, n15462;
    wire [13:0]PWM_DDS_accumulator_12__N_321;
    
    wire n15461, n15460, n15459, n15458;
    wire [24:0]count_24__N_543_adj_1406;
    wire [24:0]n52_adj_1407;
    
    wire n15457;
    wire [24:0]count2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(11[34:40])
    wire [24:0]count6;   // d:/fpga_project/lattice_diamond/piano/speaker.v(12[52:58])
    wire [24:0]n3400;
    
    wire n10946;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [24:0]n3546;
    wire [24:0]count4;   // d:/fpga_project/lattice_diamond/piano/speaker.v(12[14:20])
    wire [24:0]count5;   // d:/fpga_project/lattice_diamond/piano/speaker.v(12[33:39])
    wire [24:0]n3429;
    
    wire n17243, n17244, n17245, n18854, n18925, n16952, en_0__N_252, 
        n7_adj_849, n923, n18718, n18642, n16929, n903, n18712, 
        n879, n480, n18698, n10269, n16816, n18689, n18347, n18345, 
        clk_N_168_enable_524, n18857, n18858, n18968;
    wire [24:0]n3487;
    wire [24:0]n3458;
    wire [24:0]n3600;
    
    wire n12287, n18732, n18818, n18764, n18970, n18967, clk_N_168_enable_523, 
        n18817, n18665, n18662, n4, n17;
    wire [24:0]n2682;
    wire [24:0]n2713;
    
    wire n3082;
    wire [24:0]n2779;
    
    wire n18966, n17242, n10879;
    wire [24:0]count13;   // d:/fpga_project/lattice_diamond/piano/speaker.v(15[14:21])
    wire [24:0]n3573;
    wire [24:0]u_count2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[33:41])
    
    wire n10964;
    wire [24:0]n3681;
    wire [17:0]cycle_17__N_740;
    
    wire n17920;
    wire [24:0]n2809;
    
    wire n18656;
    wire [24:0]n2744;
    wire [24:0]n2651;
    
    wire n3084, n14_adj_855, n3_adj_858, n17236, n17134, n18920, 
        n18664, n18762, n18919, n18653, n18675, n468;
    wire [24:0]n184;
    wire [15:0]fcw_r_adj_1408;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [24:0]n132;
    wire [24:0]n105;
    wire [24:0]n2479;
    wire [24:0]n2508;
    
    wire n3076, n8;
    wire [3:0]n3796;
    
    wire n17133, n16843, n10301, n18767, n3074;
    wire [24:0]n105_adj_1409;
    wire [24:0]n132_adj_1410;
    wire [24:0]count11;   // d:/fpga_project/lattice_diamond/piano/speaker.v(14[34:41])
    wire [24:0]count7;   // d:/fpga_project/lattice_diamond/piano/speaker.v(13[14:20])
    wire [24:0]n184_adj_1411;
    wire [15:0]fcw_r_adj_1412;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n18346, n137_adj_912, n18856, n18344, n121_adj_915, n16871, 
        n18699, n18693;
    wire [24:0]n105_adj_1413;
    wire [24:0]n132_adj_1414;
    wire [24:0]n184_adj_1415;
    wire [24:0]n184_adj_1416;
    wire [15:0]fcw_r_adj_1417;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [24:0]n132_adj_1418;
    wire [24:0]n105_adj_1419;
    wire [24:0]n105_adj_1420;
    wire [24:0]n132_adj_1421;
    wire [24:0]n184_adj_1422;
    wire [24:0]n2537;
    wire [24:0]n2566;
    
    wire n3078, n18821, n18820, n18824, n18823;
    wire [24:0]count8;   // d:/fpga_project/lattice_diamond/piano/speaker.v(13[33:39])
    wire [24:0]count9;   // d:/fpga_project/lattice_diamond/piano/speaker.v(13[52:58])
    wire [1:0]en;   // d:/fpga_project/lattice_diamond/piano/speaker.v(17[12:14])
    
    wire n18827, n18826, n18830, n18829, n18659, n18833, n163, 
        n18969, n18832;
    wire [3:0]n3920;
    
    wire n18923, n18922, n18924, n18921, n16_adj_1086, n3062;
    wire [24:0]count12;   // d:/fpga_project/lattice_diamond/piano/speaker.v(14[54:61])
    wire [24:0]count10;   // d:/fpga_project/lattice_diamond/piano/speaker.v(14[14:21])
    wire [24:0]n3516;
    
    wire n16004, n3080, n3072;
    wire [24:0]n2624;
    
    wire n3070;
    wire [24:0]n2595;
    
    wire n18611, n23_adj_1092, n3068, n3066;
    wire [17:0]n358;
    wire [24:0]n3627;
    wire [24:0]n3654;
    
    wire n4_adj_1099, n15482;
    wire [3:0]n3905;
    
    wire n15925, n3599, n18663, n16899, n18661, n3064, n18660, 
        n18666, n17241, n17240;
    wire [24:0]count_24__N_543_adj_1423;
    wire [24:0]n52_adj_1424;
    wire [15:0]fcw_r_adj_1425;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15481, n15480;
    wire [3:0]n3890;
    
    wire n15479;
    wire [15:0]fcw_r_adj_1426;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [15:0]fcw_r_adj_1427;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [24:0]n52_adj_1428;
    wire [24:0]count_24__N_543_adj_1429;
    
    wire n18855;
    wire [24:0]count_24__N_543_adj_1430;
    wire [24:0]n52_adj_1431;
    wire [15:0]fcw_r_adj_1432;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n18705, n19840;
    wire [15:0]fcw_r_adj_1433;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [15:0]fcw_r_adj_1434;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n18634;
    wire [15:0]fcw_r_15__N_495;
    
    wire n16936, n15966;
    wire [7:0]n7919;
    
    wire n18716, n18608;
    
    CCU2D add_2219_4 (.A0(data_out1[2]), .B0(data_out2[2]), .C0(GND_net), 
          .D0(GND_net), .A1(data_out1[3]), .B1(data_out2[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15477), .COUT(n15478), .S0(\PWM_in_12__N_452[2] ), 
          .S1(\PWM_in_12__N_452[3] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_4.INIT0 = 16'h5666;
    defparam add_2219_4.INIT1 = 16'h5666;
    defparam add_2219_4.INJECT1_0 = "NO";
    defparam add_2219_4.INJECT1_1 = "NO";
    CCU2D add_2219_2 (.A0(\data_out1[0] ), .B0(\data_out2[0] ), .C0(GND_net), 
          .D0(GND_net), .A1(data_out1[1]), .B1(data_out2[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15477), .S1(\PWM_in_12__N_452[1] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_2.INIT0 = 16'h7000;
    defparam add_2219_2.INIT1 = 16'h5666;
    defparam add_2219_2.INJECT1_0 = "NO";
    defparam add_2219_2.INJECT1_1 = "NO";
    FD1S1I rom1_4__I_6_i1 (.D(\rom1_4__N_338[0] ), .CK(rom1_4__N_289), .CD(n9292), 
           .Q(rom1[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(255[1] 306[5])
    defparam rom1_4__I_6_i1.GSR = "DISABLED";
    FD1S1I rom2_4__I_7_i1 (.D(rom2_4__N_397[0]), .CK(rom2_4__N_297), .CD(n9292), 
           .Q(\rom2[0] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam rom2_4__I_7_i1.GSR = "DISABLED";
    FD1S3AX u_count1_i1 (.D(u_count1_24__N_142[14]), .CK(clk_N_168), .Q(u_count1[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i1.GSR = "DISABLED";
    LUT4 i7746_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[21]), .C(\key_value[4] ), 
         .Z(n52[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7746_2_lut_3_lut_3_lut.init = 16'h8c8c;
    FD1S3DX PWM_DDS_accumulator_i0 (.D(n4943[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_DDS_accumulator[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i0.GSR = "DISABLED";
    FD1S3DX PWM_in__i0 (.D(n28[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i0.GSR = "DISABLED";
    FD1P3AY yinjie_box_i0 (.D(\yinjie_box_2__N_394[0] ), .SP(stat), .CK(clk_N_168), 
            .Q(fcw_r_15__N_527[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(356[8] 368[5])
    defparam yinjie_box_i0.GSR = "DISABLED";
    FD1P3AX yinjie_box_i1 (.D(\yinjie_box_2__N_394[1] ), .SP(stat), .CK(clk_N_168), 
            .Q(yinjie_box[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(356[8] 368[5])
    defparam yinjie_box_i1.GSR = "DISABLED";
    LUT4 i7609_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[7]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7609_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7610_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[8]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7610_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX i12624 (.BLUT(n18851), .ALUT(n18852), .C0(n19846), .Z(n3086));
    PFUMX i12600 (.BLUT(n18598), .ALUT(n18597), .C0(\rom2[0] ), .Z(n18599));
    FD1S1I rom1_4__I_6_i2 (.D(n3836[1]), .CK(rom1_4__N_289), .CD(n18644), 
           .Q(rom1[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(255[1] 306[5])
    defparam rom1_4__I_6_i2.GSR = "DISABLED";
    FD1S1I rom1_4__I_6_i3 (.D(n16818), .CK(rom1_4__N_289), .CD(n18622), 
           .Q(rom1[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(255[1] 306[5])
    defparam rom1_4__I_6_i3.GSR = "DISABLED";
    FD1S1I rom1_4__I_6_i4 (.D(n15957), .CK(rom1_4__N_289), .CD(n16916), 
           .Q(rom1[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(255[1] 306[5])
    defparam rom1_4__I_6_i4.GSR = "DISABLED";
    FD1S1I rom2_4__I_7_i2 (.D(n16903), .CK(rom2_4__N_297), .CD(n18643), 
           .Q(\rom2[1] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam rom2_4__I_7_i2.GSR = "DISABLED";
    FD1S1I rom2_4__I_7_i3 (.D(n16823), .CK(rom2_4__N_297), .CD(n18621), 
           .Q(rom2[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam rom2_4__I_7_i3.GSR = "DISABLED";
    FD1S1I rom2_4__I_7_i4 (.D(n15938), .CK(rom2_4__N_297), .CD(n16930), 
           .Q(\rom2[3] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam rom2_4__I_7_i4.GSR = "DISABLED";
    LUT4 i7740_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[15]), .C(\key_value[4] ), 
         .Z(n52[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7740_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7723_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[23]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7723_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7786_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[24]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7786_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i11_3_lut (.A(count1[24]), .B(count3[24]), .C(\rom2[1] ), 
         .Z(n3371[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i11_3_lut.init = 16'hcaca;
    PFUMX i12596 (.BLUT(n18592), .ALUT(n18591), .C0(\rom2[1] ), .Z(n17004));
    LUT4 i7710_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[10]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7710_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7711_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[11]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7711_2_lut_3_lut_3_lut.init = 16'h8c8c;
    CCU2D add_2216_14 (.A0(PWM_DDS_accumulator[12]), .B0(PWM_in[12]), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15462), .S0(PWM_DDS_accumulator_12__N_321[12]), .S1(PWM_DDS_accumulator_12__N_321[13]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_14.INIT0 = 16'h5666;
    defparam add_2216_14.INIT1 = 16'h0000;
    defparam add_2216_14.INJECT1_0 = "NO";
    defparam add_2216_14.INJECT1_1 = "NO";
    CCU2D add_2216_12 (.A0(PWM_DDS_accumulator[10]), .B0(PWM_in[10]), .C0(GND_net), 
          .D0(GND_net), .A1(PWM_DDS_accumulator[11]), .B1(PWM_in[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n15461), .COUT(n15462), .S0(PWM_DDS_accumulator_12__N_321[10]), 
          .S1(PWM_DDS_accumulator_12__N_321[11]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_12.INIT0 = 16'h5666;
    defparam add_2216_12.INIT1 = 16'h5666;
    defparam add_2216_12.INJECT1_0 = "NO";
    defparam add_2216_12.INJECT1_1 = "NO";
    CCU2D add_2216_10 (.A0(PWM_DDS_accumulator[8]), .B0(PWM_in[8]), .C0(GND_net), 
          .D0(GND_net), .A1(PWM_DDS_accumulator[9]), .B1(PWM_in[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15460), .COUT(n15461), .S0(PWM_DDS_accumulator_12__N_321[8]), 
          .S1(PWM_DDS_accumulator_12__N_321[9]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_10.INIT0 = 16'h5666;
    defparam add_2216_10.INIT1 = 16'h5666;
    defparam add_2216_10.INJECT1_0 = "NO";
    defparam add_2216_10.INJECT1_1 = "NO";
    CCU2D add_2216_8 (.A0(PWM_DDS_accumulator[6]), .B0(PWM_in[6]), .C0(GND_net), 
          .D0(GND_net), .A1(PWM_DDS_accumulator[7]), .B1(PWM_in[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15459), .COUT(n15460), .S0(PWM_DDS_accumulator_12__N_321[6]), 
          .S1(PWM_DDS_accumulator_12__N_321[7]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_8.INIT0 = 16'h5666;
    defparam add_2216_8.INIT1 = 16'h5666;
    defparam add_2216_8.INJECT1_0 = "NO";
    defparam add_2216_8.INJECT1_1 = "NO";
    CCU2D add_2216_6 (.A0(PWM_DDS_accumulator[4]), .B0(PWM_in[4]), .C0(GND_net), 
          .D0(GND_net), .A1(PWM_DDS_accumulator[5]), .B1(PWM_in[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15458), .COUT(n15459), .S0(PWM_DDS_accumulator_12__N_321[4]), 
          .S1(PWM_DDS_accumulator_12__N_321[5]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_6.INIT0 = 16'h5666;
    defparam add_2216_6.INIT1 = 16'h5666;
    defparam add_2216_6.INJECT1_0 = "NO";
    defparam add_2216_6.INJECT1_1 = "NO";
    LUT4 i7584_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[7]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7584_2_lut_3_lut_3_lut.init = 16'h8c8c;
    CCU2D add_2216_4 (.A0(PWM_DDS_accumulator[2]), .B0(PWM_in[2]), .C0(GND_net), 
          .D0(GND_net), .A1(PWM_DDS_accumulator[3]), .B1(PWM_in[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15457), .COUT(n15458), .S0(PWM_DDS_accumulator_12__N_321[2]), 
          .S1(PWM_DDS_accumulator_12__N_321[3]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_4.INIT0 = 16'h5666;
    defparam add_2216_4.INIT1 = 16'h5666;
    defparam add_2216_4.INJECT1_0 = "NO";
    defparam add_2216_4.INJECT1_1 = "NO";
    CCU2D add_2216_2 (.A0(PWM_DDS_accumulator[0]), .B0(PWM_in[0]), .C0(GND_net), 
          .D0(GND_net), .A1(PWM_DDS_accumulator[1]), .B1(PWM_in[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15457), .S1(PWM_DDS_accumulator_12__N_321[1]));   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[29:63])
    defparam add_2216_2.INIT0 = 16'h7000;
    defparam add_2216_2.INIT1 = 16'h5666;
    defparam add_2216_2.INJECT1_0 = "NO";
    defparam add_2216_2.INJECT1_1 = "NO";
    LUT4 mux_1603_i10_3_lut (.A(count2[23]), .B(count6[23]), .C(rom2[2]), 
         .Z(n3400[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i10_3_lut.init = 16'hcaca;
    LUT4 i7749_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[24]), .C(\key_value[4] ), 
         .Z(n52[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7749_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i7_3_lut (.A(count1[20]), .B(count3[20]), .C(\rom2[1] ), 
         .Z(n3371[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i7_3_lut.init = 16'hcaca;
    LUT4 i6021_3_lut (.A(\key_value[11] ), .B(\key_value[12] ), .C(\rom2[0] ), 
         .Z(n10946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(373[3] 428[17])
    defparam i6021_3_lut.init = 16'hcaca;
    LUT4 i7767_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[5]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7767_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7747_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[22]), .C(\key_value[4] ), 
         .Z(n52[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7747_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1603_i11_3_lut (.A(count2[24]), .B(count6[24]), .C(rom2[2]), 
         .Z(n3400[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i11_3_lut.init = 16'hcaca;
    LUT4 i7763_3_lut_4_lut_4_lut (.A(n19846), .B(count2[1]), .C(fcw_r[6]), 
         .D(\key_value[1] ), .Z(n52_adj_1405[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7763_3_lut_4_lut_4_lut.init = 16'h283c;
    FD1S3AX u_count1_i11 (.D(u_count1_24__N_142[24]), .CK(clk_N_168), .Q(u_count1[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i11.GSR = "DISABLED";
    FD1S3AX u_count1_i10 (.D(u_count1_24__N_142[23]), .CK(clk_N_168), .Q(u_count1[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i10.GSR = "DISABLED";
    FD1S3AX u_count1_i9 (.D(u_count1_24__N_142[22]), .CK(clk_N_168), .Q(u_count1[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i9.GSR = "DISABLED";
    FD1S3AX u_count1_i8 (.D(u_count1_24__N_142[21]), .CK(clk_N_168), .Q(u_count1[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i8.GSR = "DISABLED";
    FD1S3AX u_count1_i7 (.D(u_count1_24__N_142[20]), .CK(clk_N_168), .Q(u_count1[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i7.GSR = "DISABLED";
    FD1S3AX u_count1_i6 (.D(u_count1_24__N_142[19]), .CK(clk_N_168), .Q(u_count1[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i6.GSR = "DISABLED";
    FD1S3AX u_count1_i5 (.D(u_count1_24__N_142[18]), .CK(clk_N_168), .Q(u_count1[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i5.GSR = "DISABLED";
    LUT4 i11999_3_lut (.A(n3400[14]), .B(n3371[14]), .C(\rom2[0] ), .Z(n3546[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11999_3_lut.init = 16'hcaca;
    FD1S3AX u_count1_i4 (.D(u_count1_24__N_142[17]), .CK(clk_N_168), .Q(u_count1[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i4.GSR = "DISABLED";
    FD1S3AX u_count1_i3 (.D(u_count1_24__N_142[16]), .CK(clk_N_168), .Q(u_count1[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i3.GSR = "DISABLED";
    LUT4 mux_1609_i1_3_lut (.A(count4[14]), .B(count5[14]), .C(\rom2[0] ), 
         .Z(n3429[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i1_3_lut.init = 16'hcaca;
    PFUMX i11954 (.BLUT(n17243), .ALUT(n17244), .C0(rom1[1]), .Z(n17245));
    FD1S3AX u_count1_i2 (.D(u_count1_24__N_142[15]), .CK(clk_N_168), .Q(u_count1[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(311[8] 354[5])
    defparam u_count1_i2.GSR = "DISABLED";
    LUT4 n16967_bdd_3_lut_else_3_lut (.A(\key_flag[8] ), .B(\key_flag[0] ), 
         .C(\rom2[3] ), .Z(n18854)) /* synthesis lut_function=(!(A (B+(C))+!A !((C)+!B))) */ ;
    defparam n16967_bdd_3_lut_else_3_lut.init = 16'h5353;
    LUT4 i7590_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[13]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7590_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 equal_1577_i5_2_lut (.A(rom1[0]), .B(rom1[1]), .Z(n5)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(475[53:68])
    defparam equal_1577_i5_2_lut.init = 16'hdddd;
    LUT4 mux_63_Mux_16_i7_4_lut_4_lut_4_lut (.A(n18808), .B(\note[0] ), 
         .C(\note[1] ), .D(n18737), .Z(n7)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C)))) */ ;
    defparam mux_63_Mux_16_i7_4_lut_4_lut_4_lut.init = 16'h4240;
    LUT4 n17910_bdd_2_lut_4_lut (.A(n18925), .B(n16952), .C(rom1[2]), 
         .D(n19846), .Z(en_0__N_252)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n17910_bdd_2_lut_4_lut.init = 16'hffca;
    LUT4 i7735_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[10]), .C(\key_value[4] ), 
         .Z(n52[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7735_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7773_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[11]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7773_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 n10154_bdd_4_lut_4_lut (.A(n18807), .B(n18803), .C(n18737), .D(n18808), 
         .Z(n18307)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(333[11:18])
    defparam n10154_bdd_4_lut_4_lut.init = 16'h7344;
    LUT4 i12009_3_lut (.A(n3400[24]), .B(n3371[24]), .C(\rom2[0] ), .Z(n3546[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12009_3_lut.init = 16'hcaca;
    LUT4 equal_1575_i6_2_lut (.A(rom1[2]), .B(rom1[3]), .Z(n6)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(469[53:68])
    defparam equal_1575_i6_2_lut.init = 16'hbbbb;
    LUT4 i12011_3_lut (.A(n3400[23]), .B(n3371[23]), .C(\rom2[0] ), .Z(n3546[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12011_3_lut.init = 16'hcaca;
    LUT4 mux_57_i18_4_lut_4_lut (.A(n18807), .B(n19846), .C(n7_adj_849), 
         .D(n18610), .Z(\cycle_17__N_663[17] )) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C)+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(333[11:18])
    defparam mux_57_i18_4_lut_4_lut.init = 16'h4073;
    LUT4 i12013_3_lut (.A(n3400[22]), .B(n3371[22]), .C(\rom2[0] ), .Z(n3546[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12013_3_lut.init = 16'hcaca;
    LUT4 i12015_3_lut (.A(n3400[21]), .B(n3371[21]), .C(\rom2[0] ), .Z(n3546[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12015_3_lut.init = 16'hcaca;
    LUT4 i12017_3_lut (.A(n3400[20]), .B(n3371[20]), .C(\rom2[0] ), .Z(n3546[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12017_3_lut.init = 16'hcaca;
    LUT4 i12019_3_lut (.A(n3400[19]), .B(n3371[19]), .C(\rom2[0] ), .Z(n3546[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12019_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n923), .B(n18718), .C(n18642), .D(n16929), 
         .Z(n16823)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(475[13] 479[21])
    defparam i1_3_lut_4_lut.init = 16'hff0e;
    LUT4 i12021_3_lut (.A(n3400[18]), .B(n3371[18]), .C(\rom2[0] ), .Z(n3546[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12021_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_rep_460_4_lut (.A(n18719), .B(n911), .C(n903), .D(n907), 
         .Z(n18642)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(469[13] 479[21])
    defparam i3_3_lut_rep_460_4_lut.init = 16'hfffe;
    LUT4 i12023_3_lut (.A(n3400[17]), .B(n3371[17]), .C(\rom2[0] ), .Z(n3546[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12023_3_lut.init = 16'hcaca;
    LUT4 i12025_3_lut (.A(n3400[16]), .B(n3371[16]), .C(\rom2[0] ), .Z(n3546[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12025_3_lut.init = 16'hcaca;
    LUT4 i12027_3_lut (.A(n3400[15]), .B(n3371[15]), .C(\rom2[0] ), .Z(n3546[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12027_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(n895), .B(n18677), .C(n887), .D(n891), .Z(n16929)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(457[13] 479[21])
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_rep_439_3_lut_4_lut (.A(n18712), .B(n879), .C(n9292), 
         .D(n18713), .Z(n18621)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(482[8:20])
    defparam i2_2_lut_rep_439_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut (.A(n480), .B(n18698), .C(n10269), .Z(n15957)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[13] 300[21])
    defparam i2_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_31 (.A(n480), .B(n18698), .C(n10269), .D(n16816), 
         .Z(n16818)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[13] 300[21])
    defparam i1_3_lut_4_lut_adj_31.init = 16'hff0e;
    LUT4 i2_3_lut_4_lut_adj_32 (.A(n456), .B(n18689), .C(n444), .D(n11464), 
         .Z(n16816)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(278[13] 300[21])
    defparam i2_3_lut_4_lut_adj_32.init = 16'hfffe;
    LUT4 i2_2_lut_rep_440_3_lut_4_lut (.A(n18676), .B(n436), .C(n18679), 
         .D(n9292), .Z(n18622)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[13] 300[21])
    defparam i2_2_lut_rep_440_3_lut_4_lut.init = 16'hfffe;
    LUT4 n18347_bdd_4_lut (.A(n18347), .B(n18345), .C(\rom2[0] ), .D(n19846), 
         .Z(clk_N_168_enable_524)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;
    defparam n18347_bdd_4_lut.init = 16'hff35;
    LUT4 n18857_bdd_3_lut_12887 (.A(n18857), .B(n18858), .C(rom1[3]), 
         .Z(n18968)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n18857_bdd_3_lut_12887.init = 16'h3535;
    LUT4 equal_1574_i5_2_lut (.A(rom1[0]), .B(rom1[1]), .Z(n5_adj_11)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(466[51:66])
    defparam equal_1574_i5_2_lut.init = 16'hbbbb;
    LUT4 i12040_3_lut (.A(n3487[14]), .B(n3458[14]), .C(\rom2[1] ), .Z(n3600[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12040_3_lut.init = 16'hcaca;
    LUT4 n17246_bdd_3_lut_then_3_lut (.A(\key_flag[9] ), .B(\key_flag[10] ), 
         .C(rom1[0]), .Z(n18858)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n17246_bdd_3_lut_then_3_lut.init = 16'h3535;
    LUT4 i7435_2_lut (.A(rom1[2]), .B(rom1[3]), .Z(n12287)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7435_2_lut.init = 16'h8888;
    LUT4 i18_4_lut_4_lut_then_4_lut (.A(n18732), .B(\note[4] ), .C(\note[3] ), 
         .D(\note[2] ), .Z(n18818)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C (D)+!C !(D)))+!A)) */ ;
    defparam i18_4_lut_4_lut_then_4_lut.init = 16'h2082;
    LUT4 equal_1555_i6_2_lut_rep_565 (.A(rom2[2]), .B(\rom2[3] ), .Z(n18747)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[51:65])
    defparam equal_1555_i6_2_lut_rep_565.init = 16'hdddd;
    LUT4 i105_3_lut_rep_507_4_lut (.A(rom2[2]), .B(\rom2[3] ), .C(n18764), 
         .D(n18754), .Z(n18689)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[51:65])
    defparam i105_3_lut_rep_507_4_lut.init = 16'hfd00;
    LUT4 n18971_bdd_2_lut_4_lut (.A(n18970), .B(n18967), .C(rom1[2]), 
         .D(n19846), .Z(clk_N_168_enable_523)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n18971_bdd_2_lut_4_lut.init = 16'hffca;
    LUT4 n17246_bdd_3_lut_else_3_lut (.A(\key_flag[1] ), .B(\key_flag[2] ), 
         .C(rom1[0]), .Z(n18857)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n17246_bdd_3_lut_else_3_lut.init = 16'h3535;
    LUT4 i18_4_lut_4_lut_else_4_lut (.A(rom1[2]), .B(rom1[3]), .C(rom1[0]), 
         .D(rom1[1]), .Z(n18817)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i18_4_lut_4_lut_else_4_lut.init = 16'h0100;
    LUT4 i4516_2_lut_rep_483_4_lut (.A(n18722), .B(n12156), .C(n18724), 
         .D(n436), .Z(n18665)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[16:65])
    defparam i4516_2_lut_rep_483_4_lut.init = 16'hffa2;
    LUT4 i1_2_lut_rep_480_4_lut (.A(n18720), .B(n18813), .C(n6_adj_12), 
         .D(n895), .Z(n18662)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(457[16:65])
    defparam i1_2_lut_rep_480_4_lut.init = 16'hffa2;
    LUT4 equal_1570_i6_2_lut (.A(rom1[2]), .B(rom1[3]), .Z(n6_adj_12)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(454[51:65])
    defparam equal_1570_i6_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut (.A(n18763), .B(n4), .C(n18761), .D(n16917), 
         .Z(n17)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i1_4_lut_4_lut.init = 16'h5051;
    LUT4 i7549_4_lut_4_lut (.A(n18763), .B(n9654), .C(n16909), .D(n10160), 
         .Z(n406)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i7549_4_lut_4_lut.init = 16'h5150;
    L6MUX21 mux_1501_i11 (.D0(n2682[24]), .D1(n2713[24]), .SD(n3082), 
            .Z(n2779[24]));
    L6MUX21 mux_1501_i10 (.D0(n2682[23]), .D1(n2713[23]), .SD(n3082), 
            .Z(n2779[23]));
    LUT4 i7547_4_lut_4_lut (.A(n18763), .B(n18755), .C(n18667), .D(n18761), 
         .Z(n410)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i7547_4_lut_4_lut.init = 16'h5540;
    LUT4 i7712_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[12]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7712_2_lut_3_lut_3_lut.init = 16'h8c8c;
    L6MUX21 mux_1501_i9 (.D0(n2682[22]), .D1(n2713[22]), .SD(n3082), .Z(n2779[22]));
    L6MUX21 mux_1501_i8 (.D0(n2682[21]), .D1(n2713[21]), .SD(n3082), .Z(n2779[21]));
    L6MUX21 mux_1501_i7 (.D0(n2682[20]), .D1(n2713[20]), .SD(n3082), .Z(n2779[20]));
    L6MUX21 mux_1501_i6 (.D0(n2682[19]), .D1(n2713[19]), .SD(n3082), .Z(n2779[19]));
    LUT4 n17245_bdd_3_lut_12869 (.A(n17245), .B(n18966), .C(rom1[3]), 
         .Z(n18967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n17245_bdd_3_lut_12869.init = 16'hcaca;
    L6MUX21 mux_1501_i5 (.D0(n2682[18]), .D1(n2713[18]), .SD(n3082), .Z(n2779[18]));
    L6MUX21 mux_1501_i4 (.D0(n2682[17]), .D1(n2713[17]), .SD(n3082), .Z(n2779[17]));
    LUT4 i11669_4_lut (.A(n17242), .B(rom1[1]), .C(rom1[3]), .D(n10879), 
         .Z(n16952)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B (C (D))))) */ ;
    defparam i11669_4_lut.init = 16'h0535;
    L6MUX21 mux_1501_i3 (.D0(n2682[16]), .D1(n2713[16]), .SD(n3082), .Z(n2779[16]));
    LUT4 i55_3_lut_4_lut (.A(n18755), .B(n18815), .C(n31), .D(n18720), 
         .Z(n321)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(284[16:49])
    defparam i55_3_lut_4_lut.init = 16'h1110;
    L6MUX21 mux_1501_i2 (.D0(n2682[15]), .D1(n2713[15]), .SD(n3082), .Z(n2779[15]));
    FD1S3DX PWM_in__i12 (.D(n28[12]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i12.GSR = "DISABLED";
    LUT4 equal_1566_i6_2_lut (.A(rom1[2]), .B(rom1[3]), .Z(n6_adj_13)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(442[51:65])
    defparam equal_1566_i6_2_lut.init = 16'heeee;
    LUT4 mux_1607_i8_3_lut (.A(n3429[21]), .B(count13[21]), .C(\rom2[3] ), 
         .Z(n3573[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i8_3_lut.init = 16'hcaca;
    FD1S3DX PWM_in__i11 (.D(n28[11]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i11.GSR = "DISABLED";
    FD1S3DX PWM_in__i10 (.D(n28[10]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i10.GSR = "DISABLED";
    FD1S3DX PWM_in__i9 (.D(n28[9]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i9.GSR = "DISABLED";
    FD1S3DX PWM_in__i8 (.D(n28[8]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i8.GSR = "DISABLED";
    FD1S3DX PWM_in__i7 (.D(n28[7]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i7.GSR = "DISABLED";
    FD1S3DX PWM_in__i6 (.D(n28[6]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i6.GSR = "DISABLED";
    FD1S3DX PWM_in__i5 (.D(n28[5]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i5.GSR = "DISABLED";
    FD1S3DX PWM_in__i4 (.D(n28[4]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i4.GSR = "DISABLED";
    FD1S3DX PWM_in__i3 (.D(n28[3]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i3.GSR = "DISABLED";
    FD1S3DX PWM_in__i2 (.D(n28[2]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i2.GSR = "DISABLED";
    FD1S3DX PWM_in__i1 (.D(n28[1]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(PWM_in[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(553[10] 556[22])
    defparam PWM_in__i1.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i13 (.D(PWM_DDS_accumulator_12__N_321[13]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(pwm_out2_c)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i13.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i12 (.D(PWM_DDS_accumulator_12__N_321[12]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i12.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i11 (.D(PWM_DDS_accumulator_12__N_321[11]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i11.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i10 (.D(PWM_DDS_accumulator_12__N_321[10]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i10.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i9 (.D(PWM_DDS_accumulator_12__N_321[9]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i9.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i8 (.D(PWM_DDS_accumulator_12__N_321[8]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i8.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i7 (.D(PWM_DDS_accumulator_12__N_321[7]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i7.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i6 (.D(PWM_DDS_accumulator_12__N_321[6]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i6.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i5 (.D(PWM_DDS_accumulator_12__N_321[5]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i5.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i4 (.D(PWM_DDS_accumulator_12__N_321[4]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i4.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i3 (.D(PWM_DDS_accumulator_12__N_321[3]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i3.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i2 (.D(PWM_DDS_accumulator_12__N_321[2]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i2.GSR = "DISABLED";
    FD1S3DX PWM_DDS_accumulator_i1 (.D(PWM_DDS_accumulator_12__N_321[1]), 
            .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(PWM_DDS_accumulator[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(546[6:64])
    defparam PWM_DDS_accumulator_i1.GSR = "DISABLED";
    FD1S3IX u_count2_i11 (.D(n3681[24]), .CK(clk_N_168), .CD(n10964), 
            .Q(u_count2[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i11.GSR = "DISABLED";
    PFUMX i6399 (.BLUT(n17), .ALUT(cycle_17__N_740[7]), .C0(n19846), .Z(\cycle_17__N_663[7] ));
    LUT4 n17920_bdd_2_lut (.A(n17920), .B(n19846), .Z(n10964)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n17920_bdd_2_lut.init = 16'heeee;
    FD1S3IX u_count2_i10 (.D(n3681[23]), .CK(clk_N_168), .CD(n10964), 
            .Q(u_count2[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i10.GSR = "DISABLED";
    FD1S3IX u_count2_i9 (.D(n3681[22]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i9.GSR = "DISABLED";
    FD1S3IX u_count2_i8 (.D(n3681[21]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i8.GSR = "DISABLED";
    FD1S3IX u_count2_i7 (.D(n3681[20]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i7.GSR = "DISABLED";
    FD1S3IX u_count2_i6 (.D(n3681[19]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i6.GSR = "DISABLED";
    FD1S3IX u_count2_i5 (.D(n3681[18]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i5.GSR = "DISABLED";
    FD1S3IX u_count2_i4 (.D(n3681[17]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i4.GSR = "DISABLED";
    FD1S3IX u_count2_i3 (.D(n3681[16]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i3.GSR = "DISABLED";
    FD1S3IX u_count2_i2 (.D(n3681[15]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i2.GSR = "DISABLED";
    LUT4 mux_63_Mux_12_i15_4_lut_4_lut (.A(n18808), .B(n18807), .C(n14_adj_14), 
         .D(n3), .Z(\cycle_17__N_740[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam mux_63_Mux_12_i15_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_1486_i1_3_lut (.A(n2779[14]), .B(n2809[14]), .C(n3086), .Z(u_count1_24__N_142[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i1_3_lut.init = 16'hcaca;
    LUT4 i7803_4_lut_4_lut_4_lut (.A(n18808), .B(n18656), .C(n18772), 
         .D(n18807), .Z(cycle_17__N_740[2])) /* synthesis lut_function=(!(A ((D)+!B)+!A ((D)+!C))) */ ;
    defparam i7803_4_lut_4_lut_4_lut.init = 16'h00d8;
    L6MUX21 mux_1501_i1 (.D0(n2682[14]), .D1(n2713[14]), .SD(n3082), .Z(n2779[14]));
    PFUMX mux_1492_i11 (.BLUT(n2744[24]), .ALUT(n2651[24]), .C0(n3084), 
          .Z(n2809[24]));
    LUT4 mux_63_Mux_11_i15_4_lut_4_lut (.A(n18808), .B(n18807), .C(n14_adj_855), 
         .D(n3_adj_15), .Z(\cycle_17__N_740[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;
    defparam mux_63_Mux_11_i15_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_63_Mux_13_i7_3_lut_4_lut_4_lut_4_lut (.A(n18808), .B(\note[1] ), 
         .C(n18737), .D(\note[0] ), .Z(n7_adj_16)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (D)) */ ;
    defparam mux_63_Mux_13_i7_3_lut_4_lut_4_lut_4_lut.init = 16'hdda8;
    LUT4 i7806_4_lut_4_lut_4_lut (.A(n18808), .B(n3_adj_858), .C(n18734), 
         .D(n18807), .Z(cycle_17__N_740[7])) /* synthesis lut_function=(!(A ((D)+!B)+!A ((D)+!C))) */ ;
    defparam i7806_4_lut_4_lut_4_lut.init = 16'h00d8;
    PFUMX mux_1492_i10 (.BLUT(n2744[23]), .ALUT(n2651[23]), .C0(n3084), 
          .Z(n2809[23]));
    LUT4 rom2_3__bdd_4_lut (.A(\rom2[3] ), .B(\rom2[0] ), .C(\rom2[1] ), 
         .D(rom2[2]), .Z(n17920)) /* synthesis lut_function=(A (C (D))+!A !(B+(C+(D)))) */ ;
    defparam rom2_3__bdd_4_lut.init = 16'ha001;
    PFUMX mux_1492_i9 (.BLUT(n2744[22]), .ALUT(n2651[22]), .C0(n3084), 
          .Z(n2809[22]));
    LUT4 i11843_3_lut (.A(n17236), .B(n10946), .C(rom2[2]), .Z(n17134)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i11843_3_lut.init = 16'h3a3a;
    PFUMX mux_1492_i8 (.BLUT(n2744[21]), .ALUT(n2651[21]), .C0(n3084), 
          .Z(n2809[21]));
    LUT4 i7771_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[9]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7771_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 key_value_7__bdd_3_lut_12872 (.A(\key_value[7] ), .B(rom1[1]), 
         .C(\key_value[9] ), .Z(n18920)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)))) */ ;
    defparam key_value_7__bdd_3_lut_12872.init = 16'h1d1d;
    PFUMX mux_1492_i7 (.BLUT(n2744[20]), .ALUT(n2651[20]), .C0(n3084), 
          .Z(n2809[20]));
    LUT4 i12083_3_lut (.A(n3487[15]), .B(n3458[15]), .C(\rom2[1] ), .Z(n3600[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12083_3_lut.init = 16'hcaca;
    LUT4 i12085_3_lut (.A(n3487[16]), .B(n3458[16]), .C(\rom2[1] ), .Z(n3600[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12085_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_482_4_lut (.A(n18754), .B(n18764), .C(n18747), .D(n456), 
         .Z(n18664)) /* synthesis lut_function=(A (B+(C+(D)))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(275[16:65])
    defparam i1_2_lut_rep_482_4_lut.init = 16'hffa8;
    LUT4 i1_2_lut_rep_576 (.A(\rom2[0] ), .B(\rom2[1] ), .Z(n18758)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam i1_2_lut_rep_576.init = 16'heeee;
    LUT4 i12087_3_lut (.A(n3487[17]), .B(n3458[17]), .C(\rom2[1] ), .Z(n3600[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12087_3_lut.init = 16'hcaca;
    LUT4 i129_3_lut_rep_516_4_lut (.A(\rom2[0] ), .B(\rom2[1] ), .C(n18762), 
         .D(n18761), .Z(n18698)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam i129_3_lut_rep_516_4_lut.init = 16'hef00;
    LUT4 i12089_3_lut (.A(n3487[18]), .B(n3458[18]), .C(\rom2[1] ), .Z(n3600[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12089_3_lut.init = 16'hcaca;
    PFUMX mux_1492_i6 (.BLUT(n2744[19]), .ALUT(n2651[19]), .C0(n3084), 
          .Z(n2809[19]));
    LUT4 i12091_3_lut (.A(n3487[19]), .B(n3458[19]), .C(\rom2[1] ), .Z(n3600[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12091_3_lut.init = 16'hcaca;
    LUT4 key_value_7__bdd_3_lut_12635 (.A(rom1[1]), .B(\key_value[8] ), 
         .C(\key_value[10] ), .Z(n18919)) /* synthesis lut_function=(!(A (C)+!A (B))) */ ;
    defparam key_value_7__bdd_3_lut_12635.init = 16'h1b1b;
    PFUMX mux_1492_i5 (.BLUT(n2744[18]), .ALUT(n2651[18]), .C0(n3084), 
          .Z(n2809[18]));
    LUT4 i10524_2_lut (.A(PWM_DDS_accumulator[0]), .B(PWM_in[0]), .Z(n4943[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i10524_2_lut.init = 16'h6666;
    LUT4 i12093_3_lut (.A(n3487[20]), .B(n3458[20]), .C(\rom2[1] ), .Z(n3600[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12093_3_lut.init = 16'hcaca;
    LUT4 i127_2_lut_rep_579 (.A(\key_value[11] ), .B(\key_flag[11] ), .Z(n18761)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(293[16:51])
    defparam i127_2_lut_rep_579.init = 16'h4444;
    LUT4 i5_2_lut_rep_471_3_lut_4_lut (.A(\key_value[11] ), .B(\key_flag[11] ), 
         .C(n18771), .D(n18763), .Z(n18653)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(293[16:51])
    defparam i5_2_lut_rep_471_3_lut_4_lut.init = 16'hfff4;
    LUT4 i317_3_lut_rep_536_4_lut (.A(\key_value[11] ), .B(\key_flag[11] ), 
         .C(n12287), .D(n18814), .Z(n18718)) /* synthesis lut_function=(!(A+!(B ((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(293[16:51])
    defparam i317_3_lut_rep_536_4_lut.init = 16'h4404;
    LUT4 i12095_3_lut (.A(n3487[21]), .B(n3458[21]), .C(\rom2[1] ), .Z(n3600[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12095_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_438_2_lut_3_lut_3_lut_4_lut (.A(\key_value[11] ), .B(\key_flag[11] ), 
         .C(n18768), .D(n18771), .Z(n18620)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(293[16:51])
    defparam i1_2_lut_rep_438_2_lut_3_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i12097_3_lut (.A(n3487[22]), .B(n3458[22]), .C(\rom2[1] ), .Z(n3600[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12097_3_lut.init = 16'hcaca;
    LUT4 i2280_4_lut (.A(n18803), .B(\note[4] ), .C(\note[2] ), .D(\note[3] ), 
         .Z(\yinjie_box_2__N_394[1] )) /* synthesis lut_function=(A (B)+!A (B+(C (D)))) */ ;
    defparam i2280_4_lut.init = 16'hdccc;
    LUT4 i12099_3_lut (.A(n3487[23]), .B(n3458[23]), .C(\rom2[1] ), .Z(n3600[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12099_3_lut.init = 16'hcaca;
    LUT4 i7453_2_lut_rep_580 (.A(rom2[2]), .B(\rom2[3] ), .Z(n18762)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7453_2_lut_rep_580.init = 16'h8888;
    LUT4 i133_3_lut_4_lut (.A(rom2[2]), .B(\rom2[3] ), .C(n5_adj_17), 
         .D(n18763), .Z(n480)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i133_3_lut_4_lut.init = 16'hf700;
    PFUMX mux_1492_i4 (.BLUT(n2744[17]), .ALUT(n2651[17]), .C0(n3084), 
          .Z(n2809[17]));
    LUT4 i131_2_lut_rep_581 (.A(\key_value[12] ), .B(\key_flag[12] ), .Z(n18763)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i131_2_lut_rep_581.init = 16'h4444;
    LUT4 i12101_3_lut (.A(n3487[24]), .B(n3458[24]), .C(\rom2[1] ), .Z(n3600[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12101_3_lut.init = 16'hcaca;
    LUT4 i5_2_lut_rep_527_3_lut_4_lut (.A(\key_value[12] ), .B(\key_flag[12] ), 
         .C(\key_flag[11] ), .D(\key_value[11] ), .Z(n18709)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i5_2_lut_rep_527_3_lut_4_lut.init = 16'h44f4;
    PFUMX mux_1492_i3 (.BLUT(n2744[16]), .ALUT(n2651[16]), .C0(n3084), 
          .Z(n2809[16]));
    LUT4 i3_2_lut_rep_493_3_lut (.A(\key_value[12] ), .B(\key_flag[12] ), 
         .C(n19846), .Z(n18675)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i3_2_lut_rep_493_3_lut.init = 16'hf4f4;
    LUT4 i321_3_lut_4_lut (.A(\key_value[12] ), .B(\key_flag[12] ), .C(n12287), 
         .D(n5), .Z(n923)) /* synthesis lut_function=(!(A+!(B ((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i321_3_lut_4_lut.init = 16'h4404;
    PFUMX mux_1492_i2 (.BLUT(n2744[15]), .ALUT(n2651[15]), .C0(n3084), 
          .Z(n2809[15]));
    LUT4 i1_2_lut_rep_582 (.A(\rom2[1] ), .B(\rom2[0] ), .Z(n18764)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_582.init = 16'hdddd;
    LUT4 i121_3_lut_4_lut (.A(\rom2[1] ), .B(\rom2[0] ), .C(n18770), .D(n18768), 
         .Z(n468)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i121_3_lut_4_lut.init = 16'hfd00;
    LUT4 i7456_3_lut_4_lut (.A(n19846), .B(\key_value[0] ), .C(n184[0]), 
         .D(fcw_r_adj_1408[0]), .Z(n132[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D))))) */ ;
    defparam i7456_3_lut_4_lut.init = 16'h0bb0;
    LUT4 i7911_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[1]), 
         .Z(n132[1])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7911_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i11 (.BLUT(n2479[24]), .ALUT(n2508[24]), .C0(n3076), 
          .Z(n2682[24]));
    LUT4 i7912_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[2]), 
         .Z(n132[2])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7912_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7913_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[3]), 
         .Z(n132[3])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7913_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i10 (.BLUT(n2479[23]), .ALUT(n2508[23]), .C0(n3076), 
          .Z(n2682[23]));
    LUT4 i7914_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[4]), 
         .Z(n132[4])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7914_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7915_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[5]), 
         .Z(n132[5])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7915_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7916_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[6]), 
         .Z(n132[6])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7916_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7917_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[7]), 
         .Z(n132[7])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7917_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7918_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[8]), 
         .Z(n132[8])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7918_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7919_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[9]), 
         .Z(n132[9])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7919_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7920_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[10]), 
         .Z(n132[10])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7920_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n18685), .B(n18619), .C(n16876), .D(n18720), 
         .Z(clk_N_168_enable_512)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[16:49])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_1581_i9 (.BLUT(n2479[22]), .ALUT(n2508[22]), .C0(n3076), 
          .Z(n2682[22]));
    LUT4 i7921_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[11]), 
         .Z(n132[11])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7921_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i8 (.BLUT(n2479[21]), .ALUT(n2508[21]), .C0(n3076), 
          .Z(n2682[21]));
    LUT4 i7922_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[12]), 
         .Z(n132[12])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7922_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7923_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[13]), 
         .Z(n132[13])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7923_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i7 (.BLUT(n2479[20]), .ALUT(n2508[20]), .C0(n3076), 
          .Z(n2682[20]));
    LUT4 i7924_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[14]), 
         .Z(n132[14])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7924_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7925_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[15]), 
         .Z(n132[15])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7925_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i6 (.BLUT(n2479[19]), .ALUT(n2508[19]), .C0(n3076), 
          .Z(n2682[19]));
    PFUMX mux_1581_i5 (.BLUT(n2479[18]), .ALUT(n2508[18]), .C0(n3076), 
          .Z(n2682[18]));
    LUT4 i7926_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[16]), 
         .Z(n132[16])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7926_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7927_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[17]), 
         .Z(n132[17])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7927_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7928_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[18]), 
         .Z(n132[18])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7928_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7929_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[19]), 
         .Z(n132[19])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7929_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7930_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[20]), 
         .Z(n132[20])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7930_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7931_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[21]), 
         .Z(n132[21])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7931_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i4 (.BLUT(n2479[17]), .ALUT(n2508[17]), .C0(n3076), 
          .Z(n2682[17]));
    LUT4 i7932_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[22]), 
         .Z(n132[22])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7932_2_lut_3_lut.init = 16'hb0b0;
    PFUMX mux_1581_i3 (.BLUT(n2479[16]), .ALUT(n2508[16]), .C0(n3076), 
          .Z(n2682[16]));
    LUT4 i7933_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[23]), 
         .Z(n132[23])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7933_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i8075_3_lut_4_lut (.A(n18736), .B(n18735), .C(n18722), .D(n18725), 
         .Z(n247)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[16:49])
    defparam i8075_3_lut_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_3_lut_4_lut_adj_33 (.A(n18736), .B(n18735), .C(n18722), 
         .D(n18725), .Z(n8)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[16:49])
    defparam i1_2_lut_3_lut_4_lut_adj_33.init = 16'h1110;
    PFUMX mux_1581_i2 (.BLUT(n2479[15]), .ALUT(n2508[15]), .C0(n3076), 
          .Z(n2682[15]));
    PFUMX mux_1492_i1 (.BLUT(n2744[14]), .ALUT(n2651[14]), .C0(n3084), 
          .Z(n2809[14]));
    LUT4 i3_2_lut_3_lut_4_lut (.A(n18736), .B(n18735), .C(n18708), .D(n18754), 
         .Z(n9)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[16:49])
    defparam i3_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i8054_4_lut_4_lut_4_lut (.A(n18768), .B(n331), .C(n18771), .D(n18709), 
         .Z(n415)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(287[16:49])
    defparam i8054_4_lut_4_lut_4_lut.init = 16'h00f4;
    LUT4 i7934_2_lut_3_lut (.A(n19846), .B(\key_value[0] ), .C(n105[24]), 
         .Z(n132[24])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7934_2_lut_3_lut.init = 16'hb0b0;
    LUT4 mux_1603_i7_3_lut (.A(count2[20]), .B(count6[20]), .C(rom2[2]), 
         .Z(n3400[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i7_3_lut.init = 16'hcaca;
    LUT4 i7724_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[24]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7724_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7502_2_lut_4_lut (.A(n18771), .B(n12156), .C(n18770), .D(n468), 
         .Z(n3796[1])) /* synthesis lut_function=(A ((C+(D))+!B)+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(290[16:68])
    defparam i7502_2_lut_4_lut.init = 16'hffa2;
    LUT4 n10154_bdd_3_lut_4_lut (.A(n18620), .B(n18755), .C(n18763), .D(n18651), 
         .Z(n18308)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+(D))))) */ ;
    defparam n10154_bdd_3_lut_4_lut.init = 16'h0e0f;
    LUT4 i12134_3_lut (.A(n18850), .B(n18599), .C(rom2[2]), .Z(n17133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i12134_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_34 (.A(rom1[0]), .B(rom1[3]), .C(rom1[1]), 
         .D(rom1[2]), .Z(n16843)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_34.init = 16'h0040;
    PFUMX mux_1581_i1 (.BLUT(n2479[14]), .ALUT(n2508[14]), .C0(n3076), 
          .Z(n2682[14]));
    LUT4 n17245_bdd_4_lut_12868 (.A(\key_flag[12] ), .B(rom1[1]), .C(\key_flag[11] ), 
         .D(rom1[0]), .Z(n18966)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam n17245_bdd_4_lut_12868.init = 16'heefc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_35 (.A(rom1[2]), .B(rom1[1]), .C(rom1[3]), 
         .D(rom1[0]), .Z(n10301)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_35.init = 16'h0002;
    LUT4 i2_3_lut_3_lut_4_lut (.A(rom1[2]), .B(rom1[1]), .C(n18767), .D(n19846), 
         .Z(n3074)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_585 (.A(rom1[0]), .B(rom1[3]), .Z(n18767)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_585.init = 16'h8888;
    LUT4 i7897_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[11]), 
         .Z(n132_adj_1410[11])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7897_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7896_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[10]), 
         .Z(n132_adj_1410[10])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7896_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7895_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[9]), 
         .Z(n132_adj_1410[9])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7895_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7894_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[8]), 
         .Z(n132_adj_1410[8])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7894_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7893_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[7]), 
         .Z(n132_adj_1410[7])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7893_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7892_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[6]), 
         .Z(n132_adj_1410[6])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7892_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7891_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[5]), 
         .Z(n132_adj_1410[5])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7891_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7890_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[4]), 
         .Z(n132_adj_1410[4])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7890_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7889_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[3]), 
         .Z(n132_adj_1410[3])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7889_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_1608_i8_3_lut (.A(count11[21]), .B(count7[21]), .C(rom2[2]), 
         .Z(n3458[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i8_3_lut.init = 16'hcaca;
    LUT4 i7888_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[2]), 
         .Z(n132_adj_1410[2])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7888_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7887_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[1]), 
         .Z(n132_adj_1410[1])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7887_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7450_3_lut_4_lut (.A(\key_value[2] ), .B(n19846), .C(n184_adj_1411[0]), 
         .D(fcw_r_adj_1412[0]), .Z(n132_adj_1410[0])) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7450_3_lut_4_lut.init = 16'h0dd0;
    LUT4 i7898_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[12]), 
         .Z(n132_adj_1410[12])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7898_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7899_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[13]), 
         .Z(n132_adj_1410[13])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7899_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7900_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[14]), 
         .Z(n132_adj_1410[14])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7900_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7901_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[15]), 
         .Z(n132_adj_1410[15])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7901_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7902_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[16]), 
         .Z(n132_adj_1410[16])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7902_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7903_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[17]), 
         .Z(n132_adj_1410[17])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7903_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7904_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[18]), 
         .Z(n132_adj_1410[18])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7904_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7905_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[19]), 
         .Z(n132_adj_1410[19])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7905_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7906_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[20]), 
         .Z(n132_adj_1410[20])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7906_2_lut_3_lut.init = 16'hd0d0;
    LUT4 n18346_bdd_3_lut (.A(n18346), .B(n17004), .C(\rom2[3] ), .Z(n18347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n18346_bdd_3_lut.init = 16'hcaca;
    LUT4 i7907_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[21]), 
         .Z(n132_adj_1410[21])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7907_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7908_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[22]), 
         .Z(n132_adj_1410[22])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7908_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7909_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[23]), 
         .Z(n132_adj_1410[23])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7909_2_lut_3_lut.init = 16'hd0d0;
    LUT4 n17004_bdd_4_lut (.A(n137_adj_912), .B(rom2[2]), .C(\key_flag[1] ), 
         .D(\rom2[1] ), .Z(n18346)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B+!(C+!(D))))) */ ;
    defparam n17004_bdd_4_lut.init = 16'h4744;
    LUT4 i7910_2_lut_3_lut (.A(\key_value[2] ), .B(n19846), .C(n105_adj_1409[24]), 
         .Z(n132_adj_1410[24])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(72[14:33])
    defparam i7910_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7782_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[20]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7782_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1608_i2_3_lut (.A(count11[15]), .B(count7[15]), .C(rom2[2]), 
         .Z(n3458[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i2_3_lut.init = 16'hcaca;
    LUT4 n17008_bdd_3_lut (.A(n18856), .B(n18344), .C(\rom2[1] ), .Z(n18345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n17008_bdd_3_lut.init = 16'hcaca;
    LUT4 n17008_bdd_4_lut (.A(n121_adj_915), .B(rom2[2]), .C(\rom2[3] ), 
         .D(\key_flag[2] ), .Z(n18344)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;
    defparam n17008_bdd_4_lut.init = 16'haaab;
    LUT4 i1_2_lut_3_lut_4_lut_adj_36 (.A(rom1[0]), .B(rom1[1]), .C(rom1[2]), 
         .D(rom1[3]), .Z(n16871)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (((D)+!C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_36.init = 16'h0060;
    LUT4 equal_1562_i6_2_lut_rep_588 (.A(rom2[2]), .B(\rom2[3] ), .Z(n18770)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(290[53:68])
    defparam equal_1562_i6_2_lut_rep_588.init = 16'hbbbb;
    LUT4 i125_3_lut_rep_517_4_lut (.A(rom2[2]), .B(\rom2[3] ), .C(n12156), 
         .D(n18771), .Z(n18699)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B !(D))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(290[53:68])
    defparam i125_3_lut_rep_517_4_lut.init = 16'hbf00;
    LUT4 equal_1559_i7_2_lut_rep_511_3_lut_4_lut (.A(rom2[2]), .B(\rom2[3] ), 
         .C(\rom2[1] ), .D(\rom2[0] ), .Z(n18693)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(290[53:68])
    defparam equal_1559_i7_2_lut_rep_511_3_lut_4_lut.init = 16'hfffb;
    LUT4 i7873_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[11]), 
         .Z(n132_adj_1414[11])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7873_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7872_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[10]), 
         .Z(n132_adj_1414[10])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7872_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7871_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[9]), 
         .Z(n132_adj_1414[9])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7871_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7870_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[8]), 
         .Z(n132_adj_1414[8])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7870_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7869_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[7]), 
         .Z(n132_adj_1414[7])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7869_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7868_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[6]), 
         .Z(n132_adj_1414[6])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7868_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7783_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[21]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7783_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7867_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[5]), 
         .Z(n132_adj_1414[5])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7867_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7866_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[4]), 
         .Z(n132_adj_1414[4])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7866_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7784_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[22]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7784_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7785_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[23]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7785_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7865_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[3]), 
         .Z(n132_adj_1414[3])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7865_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7864_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[2]), 
         .Z(n132_adj_1414[2])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7864_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7863_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[1]), 
         .Z(n132_adj_1414[1])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7863_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7446_3_lut_4_lut (.A(\key_value[3] ), .B(n19846), .C(n184_adj_1415[0]), 
         .D(fcw_r_adj_1412[0]), .Z(n132_adj_1414[0])) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7446_3_lut_4_lut.init = 16'h0dd0;
    LUT4 i7874_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[12]), 
         .Z(n132_adj_1414[12])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7874_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7875_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[13]), 
         .Z(n132_adj_1414[13])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7875_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7876_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[14]), 
         .Z(n132_adj_1414[14])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7876_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7877_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[15]), 
         .Z(n132_adj_1414[15])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7877_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7878_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[16]), 
         .Z(n132_adj_1414[16])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7878_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7879_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[17]), 
         .Z(n132_adj_1414[17])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7879_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7880_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[18]), 
         .Z(n132_adj_1414[18])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7880_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7881_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[19]), 
         .Z(n132_adj_1414[19])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7881_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7882_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[20]), 
         .Z(n132_adj_1414[20])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7882_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7883_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[21]), 
         .Z(n132_adj_1414[21])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7883_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7884_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[22]), 
         .Z(n132_adj_1414[22])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7884_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7885_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[23]), 
         .Z(n132_adj_1414[23])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7885_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7886_2_lut_3_lut (.A(\key_value[3] ), .B(n19846), .C(n105_adj_1413[24]), 
         .Z(n132_adj_1414[24])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(83[14:33])
    defparam i7886_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7441_3_lut_4_lut (.A(n19846), .B(\key_value[6] ), .C(n184_adj_1416[0]), 
         .D(fcw_r_adj_1417[8]), .Z(n132_adj_1418[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D))))) */ ;
    defparam i7441_3_lut_4_lut.init = 16'h0bb0;
    LUT4 i7839_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[1]), 
         .Z(n132_adj_1418[1])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7839_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7840_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[2]), 
         .Z(n132_adj_1418[2])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7840_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7841_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[3]), 
         .Z(n132_adj_1418[3])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7841_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7842_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[4]), 
         .Z(n132_adj_1418[4])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7842_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7843_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[5]), 
         .Z(n132_adj_1418[5])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7843_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7844_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[6]), 
         .Z(n132_adj_1418[6])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7844_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7845_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[7]), 
         .Z(n132_adj_1418[7])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7845_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7846_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[8]), 
         .Z(n132_adj_1418[8])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7846_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7847_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[9]), 
         .Z(n132_adj_1418[9])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7847_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7848_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[10]), 
         .Z(n132_adj_1418[10])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7848_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7849_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[11]), 
         .Z(n132_adj_1418[11])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7849_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7850_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[12]), 
         .Z(n132_adj_1418[12])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7850_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7851_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[13]), 
         .Z(n132_adj_1418[13])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7851_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7852_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[14]), 
         .Z(n132_adj_1418[14])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7852_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7853_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[15]), 
         .Z(n132_adj_1418[15])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7853_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7854_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[16]), 
         .Z(n132_adj_1418[16])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7854_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7855_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[17]), 
         .Z(n132_adj_1418[17])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7855_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7856_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[18]), 
         .Z(n132_adj_1418[18])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7856_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7857_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[19]), 
         .Z(n132_adj_1418[19])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7857_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7858_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[20]), 
         .Z(n132_adj_1418[20])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7858_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7859_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[21]), 
         .Z(n132_adj_1418[21])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7859_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7860_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[22]), 
         .Z(n132_adj_1418[22])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7860_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7861_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[23]), 
         .Z(n132_adj_1418[23])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7861_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7862_2_lut_3_lut (.A(n19846), .B(\key_value[6] ), .C(n105_adj_1419[24]), 
         .Z(n132_adj_1418[24])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;
    defparam i7862_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i7589_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[12]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7589_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7825_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[11]), 
         .Z(n132_adj_1421[11])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7825_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7824_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[10]), 
         .Z(n132_adj_1421[10])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7824_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7823_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[9]), 
         .Z(n132_adj_1421[9])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7823_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7822_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[8]), 
         .Z(n132_adj_1421[8])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7822_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7821_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[7]), 
         .Z(n132_adj_1421[7])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7821_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7820_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[6]), 
         .Z(n132_adj_1421[6])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7820_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7819_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[5]), 
         .Z(n132_adj_1421[5])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7819_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7588_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[11]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7588_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7818_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[4]), 
         .Z(n132_adj_1421[4])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7818_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7817_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[3]), 
         .Z(n132_adj_1421[3])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7817_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7816_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[2]), 
         .Z(n132_adj_1421[2])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7816_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7815_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[1]), 
         .Z(n132_adj_1421[1])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7815_2_lut_3_lut.init = 16'hd0d0;
    PFUMX i6407 (.BLUT(n26_adj_18), .ALUT(cycle_17__N_740[2]), .C0(n19846), 
          .Z(\cycle_17__N_663[2] ));
    LUT4 i7427_3_lut_4_lut (.A(\key_value[11] ), .B(n19846), .C(n184_adj_1422[0]), 
         .D(fcw_r_adj_1412[0]), .Z(n132_adj_1421[0])) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7427_3_lut_4_lut.init = 16'h0dd0;
    LUT4 i7826_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[12]), 
         .Z(n132_adj_1421[12])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7826_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7827_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[13]), 
         .Z(n132_adj_1421[13])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7827_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7828_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[14]), 
         .Z(n132_adj_1421[14])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7828_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7829_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[15]), 
         .Z(n132_adj_1421[15])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7829_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7830_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[16]), 
         .Z(n132_adj_1421[16])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7830_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7831_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[17]), 
         .Z(n132_adj_1421[17])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7831_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7832_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[18]), 
         .Z(n132_adj_1421[18])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7832_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7833_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[19]), 
         .Z(n132_adj_1421[19])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7833_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7834_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[20]), 
         .Z(n132_adj_1421[20])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7834_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7835_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[21]), 
         .Z(n132_adj_1421[21])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7835_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7836_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[22]), 
         .Z(n132_adj_1421[22])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7836_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7837_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[23]), 
         .Z(n132_adj_1421[23])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7837_2_lut_3_lut.init = 16'hd0d0;
    PFUMX mux_1579_i2 (.BLUT(n2537[15]), .ALUT(n2566[15]), .C0(n3078), 
          .Z(n2713[15]));
    LUT4 i7838_2_lut_3_lut (.A(\key_value[11] ), .B(n19846), .C(n105_adj_1420[24]), 
         .Z(n132_adj_1421[24])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(171[14:34])
    defparam i7838_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i18_4_lut_4_lut_then_4_lut_adj_37 (.A(n18807), .B(n18808), .C(\note[1] ), 
         .D(\note[0] ), .Z(n18821)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i18_4_lut_4_lut_then_4_lut_adj_37.init = 16'h0008;
    LUT4 i18_4_lut_4_lut_else_4_lut_adj_38 (.A(rom1[3]), .B(rom1[0]), .C(rom1[1]), 
         .D(rom1[2]), .Z(n18820)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i18_4_lut_4_lut_else_4_lut_adj_38.init = 16'h0002;
    LUT4 i30_4_lut_4_lut_then_4_lut (.A(\note[0] ), .B(\note[1] ), .C(n18807), 
         .D(n18808), .Z(n18824)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i30_4_lut_4_lut_then_4_lut.init = 16'h0807;
    LUT4 i30_4_lut_4_lut_else_4_lut (.A(rom1[2]), .B(rom1[0]), .C(rom1[1]), 
         .D(rom1[3]), .Z(n18823)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (((D)+!C)+!B))) */ ;
    defparam i30_4_lut_4_lut_else_4_lut.init = 16'h006a;
    PFUMX mux_1579_i3 (.BLUT(n2537[16]), .ALUT(n2566[16]), .C0(n3078), 
          .Z(n2713[16]));
    LUT4 mux_1609_i2_3_lut (.A(count4[15]), .B(count5[15]), .C(\rom2[0] ), 
         .Z(n3429[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i2_3_lut.init = 16'hcaca;
    LUT4 i7587_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[10]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7587_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1610_i2_3_lut (.A(count8[15]), .B(count9[15]), .C(\rom2[0] ), 
         .Z(n3487[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_39 (.A(n18754), .B(n18735), .C(n18736), 
         .D(n18720), .Z(n10337)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(275[16:49])
    defparam i1_2_lut_3_lut_4_lut_adj_39.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_40 (.A(n18754), .B(n18735), .C(n18707), 
         .D(n18708), .Z(n10160)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(275[16:49])
    defparam i1_2_lut_3_lut_4_lut_adj_40.init = 16'hfffe;
    LUT4 i7586_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[9]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7586_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i6076_2_lut_3_lut_4_lut (.A(n18754), .B(n18735), .C(n18707), 
         .D(n18725), .Z(n269)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(275[16:49])
    defparam i6076_2_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i2_3_lut (.A(en[1]), .B(en[0]), .C(n19846), .Z(rom2_4__N_297)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    PFUMX mux_1579_i4 (.BLUT(n2537[17]), .ALUT(n2566[17]), .C0(n3078), 
          .Z(n2713[17]));
    LUT4 i40_4_lut_4_lut_then_4_lut (.A(n18807), .B(n18808), .C(\note[1] ), 
         .D(\note[0] ), .Z(n18827)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;
    defparam i40_4_lut_4_lut_then_4_lut.init = 16'h0440;
    LUT4 i40_4_lut_4_lut_else_4_lut (.A(rom1[1]), .B(rom1[0]), .C(rom1[2]), 
         .D(rom1[3]), .Z(n18826)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;
    defparam i40_4_lut_4_lut_else_4_lut.init = 16'h0006;
    LUT4 i18_4_lut_4_lut_then_4_lut_adj_41 (.A(n18807), .B(n18737), .C(n18803), 
         .D(n18808), .Z(n18830)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i18_4_lut_4_lut_then_4_lut_adj_41.init = 16'h4000;
    LUT4 i18_4_lut_4_lut_else_4_lut_adj_42 (.A(rom1[1]), .B(rom1[2]), .C(rom1[3]), 
         .D(rom1[0]), .Z(n18829)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i18_4_lut_4_lut_else_4_lut_adj_42.init = 16'h0040;
    LUT4 i24_4_lut_4_lut_then_3_lut (.A(\note[0] ), .B(\note[1] ), .C(n18659), 
         .Z(n18833)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i24_4_lut_4_lut_then_3_lut.init = 16'h8080;
    LUT4 n18857_bdd_4_lut_12888 (.A(n163), .B(\key_flag[0] ), .C(rom1[3]), 
         .D(rom1[0]), .Z(n18969)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B+(C+!(D))))) */ ;
    defparam n18857_bdd_4_lut_12888.init = 16'h5c5f;
    PFUMX mux_1579_i5 (.BLUT(n2537[18]), .ALUT(n2566[18]), .C0(n3078), 
          .Z(n2713[18]));
    PFUMX i12656 (.BLUT(n18969), .ALUT(n18968), .C0(rom1[1]), .Z(n18970));
    LUT4 i24_4_lut_4_lut_else_3_lut (.A(rom1[2]), .B(rom1[3]), .C(rom1[0]), 
         .D(rom1[1]), .Z(n18832)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;
    defparam i24_4_lut_4_lut_else_3_lut.init = 16'h4080;
    PFUMX mux_1579_i6 (.BLUT(n2537[19]), .ALUT(n2566[19]), .C0(n3078), 
          .Z(n2713[19]));
    LUT4 i7296_4_lut (.A(n3920[0]), .B(n18713), .C(n879), .D(n18712), 
         .Z(rom2_4__N_397[0])) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(442[13] 479[21])
    defparam i7296_4_lut.init = 16'hcfce;
    LUT4 key_value_1__bdd_2_lut_12877 (.A(\key_value[1] ), .B(rom1[1]), 
         .Z(n18923)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam key_value_1__bdd_2_lut_12877.init = 16'h4444;
    LUT4 key_value_1__bdd_3_lut_12876 (.A(\key_value[0] ), .B(rom1[1]), 
         .C(\key_value[2] ), .Z(n18922)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)))) */ ;
    defparam key_value_1__bdd_3_lut_12876.init = 16'h1d1d;
    PFUMX mux_1579_i7 (.BLUT(n2537[20]), .ALUT(n2566[20]), .C0(n3078), 
          .Z(n2713[20]));
    PFUMX mux_1579_i8 (.BLUT(n2537[21]), .ALUT(n2566[21]), .C0(n3078), 
          .Z(n2713[21]));
    LUT4 i7580_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[3]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7580_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7578_3_lut_4_lut_4_lut (.A(n19846), .B(count13[1]), .C(fcw_r_adj_1408[0]), 
         .D(\key_value[12] ), .Z(n52_adj_1407[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7578_3_lut_4_lut_4_lut.init = 16'h283c;
    PFUMX mux_1579_i9 (.BLUT(n2537[22]), .ALUT(n2566[22]), .C0(n3078), 
          .Z(n2713[22]));
    PFUMX mux_1579_i10 (.BLUT(n2537[23]), .ALUT(n2566[23]), .C0(n3078), 
          .Z(n2713[23]));
    PFUMX mux_1579_i11 (.BLUT(n2537[24]), .ALUT(n2566[24]), .C0(n3078), 
          .Z(n2713[24]));
    PFUMX mux_1579_i1 (.BLUT(n2537[14]), .ALUT(n2566[14]), .C0(n3078), 
          .Z(n2713[14]));
    LUT4 i7713_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[13]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7713_2_lut_3_lut_3_lut.init = 16'h8c8c;
    L6MUX21 i12640 (.D0(n18924), .D1(n18921), .SD(rom1[3]), .Z(n18925));
    LUT4 i7737_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[12]), .C(\key_value[4] ), 
         .Z(n52[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7737_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX i12612 (.BLUT(n18832), .ALUT(n18833), .C0(n19846), .Z(n3084));
    LUT4 i40_4_lut_4_lut_4_lut (.A(n19846), .B(n18808), .C(n16_adj_1086), 
         .D(n18709), .Z(n22_adj_19)) /* synthesis lut_function=(A (B)+!A !((D)+!C)) */ ;
    defparam i40_4_lut_4_lut_4_lut.init = 16'h88d8;
    PFUMX i12610 (.BLUT(n18829), .ALUT(n18830), .C0(n19846), .Z(n3062));
    LUT4 mux_1602_i7_3_lut (.A(count12[20]), .B(count10[20]), .C(\rom2[1] ), 
         .Z(n3516[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i7_3_lut.init = 16'hcaca;
    PFUMX i12608 (.BLUT(n18826), .ALUT(n18827), .C0(n19846), .Z(n3076));
    LUT4 i36_4_lut_4_lut (.A(n19846), .B(n18659), .C(n16004), .D(n18769), 
         .Z(n3080)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;
    defparam i36_4_lut_4_lut.init = 16'hd850;
    PFUMX i12638 (.BLUT(n18923), .ALUT(n18922), .C0(rom1[0]), .Z(n18924));
    PFUMX i12606 (.BLUT(n18823), .ALUT(n18824), .C0(n19846), .Z(n3082));
    LUT4 i7769_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[7]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7769_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7736_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[11]), .C(\key_value[4] ), 
         .Z(n52[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7736_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX i12636 (.BLUT(n18920), .ALUT(n18919), .C0(rom1[0]), .Z(n18921));
    LUT4 i7768_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[6]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7768_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1583_i1_3_lut (.A(count9[14]), .B(count10[14]), .C(n3072), 
         .Z(n2624[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i1_3_lut (.A(count7[14]), .B(count8[14]), .C(n3070), 
         .Z(n2595[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i1_3_lut.init = 16'hcaca;
    LUT4 i7766_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[4]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7766_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_2_lut_rep_429_3_lut_3_lut_4_lut_4_lut (.A(n18771), .B(n18685), 
         .C(n18709), .D(n18768), .Z(n18611)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_429_3_lut_3_lut_4_lut_4_lut.init = 16'hfffe;
    LUT4 rom2_3__bdd_4_lut_12390 (.A(\rom2[3] ), .B(rom2[2]), .C(\rom2[1] ), 
         .D(\rom2[0] ), .Z(n23_adj_1092)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)))) */ ;
    defparam rom2_3__bdd_4_lut_12390.init = 16'h6e06;
    LUT4 mux_1608_i1_3_lut (.A(count11[14]), .B(count7[14]), .C(rom2[2]), 
         .Z(n3458[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n18771), .B(n18675), .C(n18761), 
         .D(n18768), .Z(n16920)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_430_3_lut_3_lut_4_lut_4_lut (.A(n18771), .B(n18755), 
         .C(n18761), .D(n18768), .Z(n18612)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_430_3_lut_3_lut_4_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1582_i1_3_lut (.A(count11[14]), .B(count13[14]), .C(n3074), 
         .Z(n2651[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1585_i1_3_lut (.A(count5[14]), .B(count6[14]), .C(n3068), 
         .Z(n2566[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i1_3_lut.init = 16'hcaca;
    LUT4 i11675_2_lut_2_lut_3_lut_4_lut_4_lut (.A(n18771), .B(n18768), .C(n18815), 
         .D(n18755), .Z(n16959)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11675_2_lut_2_lut_3_lut_4_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1610_i1_3_lut (.A(count8[14]), .B(count9[14]), .C(\rom2[0] ), 
         .Z(n3487[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i1_3_lut.init = 16'hcaca;
    PFUMX i12604 (.BLUT(n18820), .ALUT(n18821), .C0(n19846), .Z(n3070));
    LUT4 mux_1588_i1_3_lut (.A(count3[14]), .B(count4[14]), .C(n3066), 
         .Z(n2537[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_441_2_lut_3_lut_4_lut_4_lut (.A(n18771), .B(n18768), 
         .C(n18708), .D(n18755), .Z(n18623)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_441_2_lut_3_lut_4_lut_4_lut.init = 16'hfffe;
    LUT4 mux_1585_i11_3_lut (.A(count5[24]), .B(count6[24]), .C(n3068), 
         .Z(n2566[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i11_3_lut (.A(count3[24]), .B(count4[24]), .C(n3066), 
         .Z(n2537[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i11_3_lut.init = 16'hcaca;
    LUT4 i12212_3_lut_4_lut_4_lut (.A(n19846), .B(n417), .C(n18808), .D(n18769), 
         .Z(\cycle_17__N_740[1] )) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam i12212_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_1585_i10_3_lut (.A(count5[23]), .B(count6[23]), .C(n3068), 
         .Z(n2566[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i10_3_lut (.A(count3[23]), .B(count4[23]), .C(n3066), 
         .Z(n2537[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1585_i9_3_lut (.A(count5[22]), .B(count6[22]), .C(n3068), 
         .Z(n2566[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i9_3_lut (.A(count3[22]), .B(count4[22]), .C(n3066), 
         .Z(n2537[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1585_i8_3_lut (.A(count5[21]), .B(count6[21]), .C(n3068), 
         .Z(n2566[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i8_3_lut (.A(count3[21]), .B(count4[21]), .C(n3066), 
         .Z(n2537[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1585_i7_3_lut (.A(count5[20]), .B(count6[20]), .C(n3068), 
         .Z(n2566[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i7_3_lut (.A(count3[20]), .B(count4[20]), .C(n3066), 
         .Z(n2537[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1585_i6_3_lut (.A(count5[19]), .B(count6[19]), .C(n3068), 
         .Z(n2566[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i6_3_lut (.A(count3[19]), .B(count4[19]), .C(n3066), 
         .Z(n2537[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i6_3_lut.init = 16'hcaca;
    LUT4 mux_63_Mux_14_i15_4_lut_4_lut (.A(n19846), .B(n18709), .C(n358[14]), 
         .D(n18697), .Z(\cycle_17__N_740[14] )) /* synthesis lut_function=(A (D)+!A (B+(C))) */ ;
    defparam mux_63_Mux_14_i15_4_lut_4_lut.init = 16'hfe54;
    LUT4 i7738_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[13]), .C(\key_value[4] ), 
         .Z(n52[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7738_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7739_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[14]), .C(\key_value[4] ), 
         .Z(n52[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7739_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1607_i2_3_lut (.A(n3429[15]), .B(count13[15]), .C(\rom2[3] ), 
         .Z(n3573[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1585_i5_3_lut (.A(count5[18]), .B(count6[18]), .C(n3068), 
         .Z(n2566[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i5_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_4_lut (.A(rom1[3]), .B(rom1[2]), .C(rom1[1]), 
         .D(rom1[0]), .Z(n16004)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0220;
    LUT4 mux_1588_i5_3_lut (.A(count3[18]), .B(count4[18]), .C(n3066), 
         .Z(n2537[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i5_3_lut.init = 16'hcaca;
    LUT4 mux_63_Mux_17_i7_3_lut_3_lut_3_lut_4_lut_3_lut (.A(\note[1] ), .B(\note[0] ), 
         .C(n18808), .Z(n7_adj_849)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;
    defparam mux_63_Mux_17_i7_3_lut_3_lut_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_1585_i4_3_lut (.A(count5[17]), .B(count6[17]), .C(n3068), 
         .Z(n2566[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i4_3_lut.init = 16'hcaca;
    LUT4 i39_3_lut_3_lut_4_lut_3_lut (.A(\note[1] ), .B(\note[0] ), .C(n18808), 
         .Z(n19_adj_20)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)))) */ ;
    defparam i39_3_lut_3_lut_4_lut_3_lut.init = 16'h6868;
    LUT4 i14_4_lut_rep_625 (.A(\note[2] ), .B(\note[4] ), .C(\note[3] ), 
         .Z(n18807)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i14_4_lut_rep_625.init = 16'h1818;
    LUT4 mux_1588_i4_3_lut (.A(count3[17]), .B(count4[17]), .C(n3066), 
         .Z(n2537[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i4_3_lut.init = 16'hcaca;
    LUT4 i12344_2_lut_4_lut (.A(\note[2] ), .B(\note[4] ), .C(\note[3] ), 
         .D(n19846), .Z(n17110)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (B (D)+!B !(C+!(D))))) */ ;
    defparam i12344_2_lut_4_lut.init = 16'h18ff;
    LUT4 i12272_2_lut (.A(n19846), .B(en[0]), .Z(rom1_4__N_289)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12272_2_lut.init = 16'h1111;
    LUT4 i7781_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[19]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7781_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7585_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[8]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7585_2_lut_3_lut_3_lut.init = 16'h8c8c;
    L6MUX21 mux_1599_i11 (.D0(n3627[24]), .D1(n3654[24]), .SD(n23_adj_1092), 
            .Z(n3681[24]));
    L6MUX21 mux_1599_i10 (.D0(n3627[23]), .D1(n3654[23]), .SD(n23_adj_1092), 
            .Z(n3681[23]));
    LUT4 i7810_2_lut_4_lut (.A(\note[2] ), .B(\note[3] ), .C(\note[4] ), 
         .D(\note[0] ), .Z(n14_adj_855)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B (D)+!B (C+(D))))) */ ;
    defparam i7810_2_lut_4_lut.init = 16'h006d;
    LUT4 i11658_2_lut_4_lut_3_lut (.A(\note[2] ), .B(\note[3] ), .C(\note[4] ), 
         .Z(n18808)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;
    defparam i11658_2_lut_4_lut_3_lut.init = 16'h6d6d;
    L6MUX21 mux_1599_i9 (.D0(n3627[22]), .D1(n3654[22]), .SD(n23_adj_1092), 
            .Z(n3681[22]));
    L6MUX21 mux_1599_i8 (.D0(n3627[21]), .D1(n3654[21]), .SD(n23_adj_1092), 
            .Z(n3681[21]));
    LUT4 i7481_2_lut_rep_515_4_lut (.A(\note[2] ), .B(\note[3] ), .C(\note[4] ), 
         .D(\note[1] ), .Z(n18697)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B (D)+!B (C+(D))))) */ ;
    defparam i7481_2_lut_rep_515_4_lut.init = 16'h006d;
    L6MUX21 mux_1599_i7 (.D0(n3627[20]), .D1(n3654[20]), .SD(n23_adj_1092), 
            .Z(n3681[20]));
    L6MUX21 mux_1599_i6 (.D0(n3627[19]), .D1(n3654[19]), .SD(n23_adj_1092), 
            .Z(n3681[19]));
    LUT4 i8129_2_lut_2_lut_4_lut (.A(\note[2] ), .B(\note[3] ), .C(\note[4] ), 
         .D(\note[0] ), .Z(n12983)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B+!(C (D)))) */ ;
    defparam i8129_2_lut_2_lut_4_lut.init = 16'h9200;
    LUT4 i1_2_lut_rep_477_4_lut_3_lut (.A(\note[2] ), .B(\note[3] ), .C(\note[4] ), 
         .Z(n18659)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;
    defparam i1_2_lut_rep_477_4_lut_3_lut.init = 16'h2424;
    LUT4 i4952_2_lut_2_lut_4_lut (.A(\note[2] ), .B(\note[3] ), .C(\note[4] ), 
         .D(\note[1] ), .Z(n9757)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (B (D)+!B (C+(D)))) */ ;
    defparam i4952_2_lut_2_lut_4_lut.init = 16'hff92;
    L6MUX21 mux_1599_i5 (.D0(n3627[18]), .D1(n3654[18]), .SD(n23_adj_1092), 
            .Z(n3681[18]));
    L6MUX21 mux_1599_i4 (.D0(n3627[17]), .D1(n3654[17]), .SD(n23_adj_1092), 
            .Z(n3681[17]));
    L6MUX21 mux_1599_i3 (.D0(n3627[16]), .D1(n3654[16]), .SD(n23_adj_1092), 
            .Z(n3681[16]));
    L6MUX21 mux_1599_i2 (.D0(n3627[15]), .D1(n3654[15]), .SD(n23_adj_1092), 
            .Z(n3681[15]));
    FD1P3AX en_0__413 (.D(en_0__N_252), .SP(clk_N_168_enable_523), .CK(clk_N_168), 
            .Q(en[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(191[8] 253[5])
    defparam en_0__413.GSR = "DISABLED";
    PFUMX i11844 (.BLUT(n17133), .ALUT(n17134), .C0(\rom2[3] ), .Z(n17135));
    LUT4 i4_2_lut_3_lut_4_lut (.A(rom1[2]), .B(rom1[1]), .C(rom1[3]), 
         .D(rom1[0]), .Z(n4_adj_1099)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i4_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i7583_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[6]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7583_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7579_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[2]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[2])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7579_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7611_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[9]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7611_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7612_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[10]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7612_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7718_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[18]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7718_2_lut_3_lut_3_lut.init = 16'h8c8c;
    CCU2D add_2219_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15482), 
          .S0(\PWM_in_12__N_452[12] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_cout.INIT0 = 16'h0000;
    defparam add_2219_cout.INIT1 = 16'h0000;
    defparam add_2219_cout.INJECT1_0 = "NO";
    defparam add_2219_cout.INJECT1_1 = "NO";
    L6MUX21 mux_1599_i1 (.D0(n3627[14]), .D1(n3654[14]), .SD(n23_adj_1092), 
            .Z(n3681[14]));
    LUT4 i7613_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[11]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7613_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1585_i3_3_lut (.A(count5[16]), .B(count6[16]), .C(n3068), 
         .Z(n2566[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i3_3_lut.init = 16'hcaca;
    LUT4 i7292_4_lut (.A(n3905[0]), .B(n887), .C(n891), .D(n895), .Z(n3920[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(451[13] 479[21])
    defparam i7292_4_lut.init = 16'h3032;
    LUT4 mux_1588_i3_3_lut (.A(count3[16]), .B(count4[16]), .C(n3066), 
         .Z(n2537[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i1_3_lut (.A(n3429[14]), .B(count13[14]), .C(\rom2[3] ), 
         .Z(n3573[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i1_3_lut.init = 16'hcaca;
    LUT4 i7614_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[12]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7614_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1585_i2_3_lut (.A(count5[15]), .B(count6[15]), .C(n3068), 
         .Z(n2566[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1585_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1588_i2_3_lut (.A(count3[15]), .B(count4[15]), .C(n3066), 
         .Z(n2537[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1588_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1609_i11_3_lut (.A(count4[24]), .B(count5[24]), .C(\rom2[0] ), 
         .Z(n3429[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1609_i10_3_lut (.A(count4[23]), .B(count5[23]), .C(\rom2[0] ), 
         .Z(n3429[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1583_i11_3_lut (.A(count9[24]), .B(count10[24]), .C(n3072), 
         .Z(n2624[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1609_i9_3_lut (.A(count4[22]), .B(count5[22]), .C(\rom2[0] ), 
         .Z(n3429[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i9_3_lut.init = 16'hcaca;
    LUT4 i8095_4_lut (.A(n444), .B(n18665), .C(n15925), .D(n11464), 
         .Z(n3836[1])) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[13] 300[21])
    defparam i8095_4_lut.init = 16'hccdc;
    LUT4 i1_4_lut (.A(n37), .B(n18664), .C(n464), .D(n3796[1]), .Z(n15925)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(278[13] 300[21])
    defparam i1_4_lut.init = 16'hcecc;
    LUT4 mux_1584_i11_3_lut (.A(count7[24]), .B(count8[24]), .C(n3070), 
         .Z(n2595[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i11_3_lut.init = 16'hcaca;
    LUT4 i7719_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[19]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7719_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1582_i11_3_lut (.A(count11[24]), .B(count13[24]), .C(n3074), 
         .Z(n2651[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i11_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(n464), .B(n3796[1]), .C(n18693), .D(n18815), .Z(n10269)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(284[13] 300[21])
    defparam i3_4_lut.init = 16'hfeee;
    LUT4 mux_1583_i10_3_lut (.A(count9[23]), .B(count10[23]), .C(n3072), 
         .Z(n2624[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i10_3_lut.init = 16'hcaca;
    PFUMX mux_1604_i11 (.BLUT(n3600[24]), .ALUT(n3573[24]), .C0(n3599), 
          .Z(n3654[24]));
    LUT4 mux_1584_i10_3_lut (.A(count7[23]), .B(count8[23]), .C(n3070), 
         .Z(n2595[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i10_3_lut (.A(count11[23]), .B(count13[23]), .C(n3074), 
         .Z(n2651[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i10_3_lut.init = 16'hcaca;
    PFUMX mux_1604_i10 (.BLUT(n3600[23]), .ALUT(n3573[23]), .C0(n3599), 
          .Z(n3654[23]));
    LUT4 mux_1583_i9_3_lut (.A(count9[22]), .B(count10[22]), .C(n3072), 
         .Z(n2624[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i9_3_lut (.A(count7[22]), .B(count8[22]), .C(n3070), 
         .Z(n2595[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i9_3_lut (.A(count11[22]), .B(count13[22]), .C(n3074), 
         .Z(n2651[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i9_3_lut.init = 16'hcaca;
    PFUMX mux_1604_i9 (.BLUT(n3600[22]), .ALUT(n3573[22]), .C0(n3599), 
          .Z(n3654[22]));
    LUT4 mux_1583_i8_3_lut (.A(count9[21]), .B(count10[21]), .C(n3072), 
         .Z(n2624[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i8_3_lut (.A(count7[21]), .B(count8[21]), .C(n3070), 
         .Z(n2595[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i8_3_lut (.A(count11[21]), .B(count13[21]), .C(n3074), 
         .Z(n2651[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1583_i7_3_lut (.A(count9[20]), .B(count10[20]), .C(n3072), 
         .Z(n2624[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i7_3_lut (.A(count7[20]), .B(count8[20]), .C(n3070), 
         .Z(n2595[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i7_3_lut (.A(count11[20]), .B(count13[20]), .C(n3074), 
         .Z(n2651[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1583_i6_3_lut (.A(count9[19]), .B(count10[19]), .C(n3072), 
         .Z(n2624[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i6_3_lut (.A(count7[19]), .B(count8[19]), .C(n3070), 
         .Z(n2595[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i6_3_lut (.A(count11[19]), .B(count13[19]), .C(n3074), 
         .Z(n2651[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i6_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_43 (.A(n887), .B(n18663), .C(n16899), .D(n891), 
         .Z(n16903)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(445[13] 479[21])
    defparam i1_4_lut_adj_43.init = 16'hccdc;
    LUT4 i1_4_lut_adj_44 (.A(n903), .B(n18662), .C(n18661), .D(n907), 
         .Z(n16899)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(457[13] 479[21])
    defparam i1_4_lut_adj_44.init = 16'hccdc;
    LUT4 i127_3_lut (.A(\key_flag[3] ), .B(\key_flag[5] ), .C(\rom2[1] ), 
         .Z(n137_adj_912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i127_3_lut.init = 16'hcaca;
    LUT4 mux_1583_i5_3_lut (.A(count9[18]), .B(count10[18]), .C(n3072), 
         .Z(n2624[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i5_3_lut (.A(count7[18]), .B(count8[18]), .C(n3070), 
         .Z(n2595[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i5_3_lut (.A(count11[18]), .B(count13[18]), .C(n3074), 
         .Z(n2651[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i5_3_lut.init = 16'hcaca;
    LUT4 i119_4_lut (.A(\key_flag[6] ), .B(\key_flag[10] ), .C(\rom2[3] ), 
         .D(rom2[2]), .Z(n121_adj_915)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i119_4_lut.init = 16'h0530;
    LUT4 mux_1583_i4_3_lut (.A(count9[17]), .B(count10[17]), .C(n3072), 
         .Z(n2624[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i4_3_lut (.A(count7[17]), .B(count8[17]), .C(n3070), 
         .Z(n2595[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i4_3_lut (.A(count11[17]), .B(count13[17]), .C(n3074), 
         .Z(n2651[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1583_i3_3_lut (.A(count9[16]), .B(count10[16]), .C(n3072), 
         .Z(n2624[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i3_3_lut (.A(count7[16]), .B(count8[16]), .C(n3070), 
         .Z(n2595[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i3_3_lut (.A(count11[16]), .B(count13[16]), .C(n3074), 
         .Z(n2651[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1583_i2_3_lut (.A(count9[15]), .B(count10[15]), .C(n3072), 
         .Z(n2624[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1583_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1584_i2_3_lut (.A(count7[15]), .B(count8[15]), .C(n3070), 
         .Z(n2595[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1584_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1582_i2_3_lut (.A(count11[15]), .B(count13[15]), .C(n3074), 
         .Z(n2651[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1582_i2_3_lut.init = 16'hcaca;
    FD1S3IX u_count2_i1 (.D(n3681[14]), .CK(clk_N_168), .CD(n10964), .Q(u_count2[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(495[8] 538[5])
    defparam u_count2_i1.GSR = "DISABLED";
    PFUMX mux_1604_i8 (.BLUT(n3600[21]), .ALUT(n3573[21]), .C0(n3599), 
          .Z(n3654[21]));
    PFUMX mux_1604_i7 (.BLUT(n3600[20]), .ALUT(n3573[20]), .C0(n3599), 
          .Z(n3654[20]));
    LUT4 i1_2_lut_rep_631 (.A(rom1[1]), .B(rom1[0]), .Z(n18813)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_631.init = 16'h8888;
    LUT4 equal_1572_i5_2_lut_rep_632 (.A(rom1[0]), .B(rom1[1]), .Z(n18814)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(460[51:65])
    defparam equal_1572_i5_2_lut_rep_632.init = 16'heeee;
    LUT4 i301_3_lut_4_lut (.A(rom1[0]), .B(rom1[1]), .C(n6), .D(n18815), 
         .Z(n903)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(460[51:65])
    defparam i301_3_lut_4_lut.init = 16'hfe00;
    LUT4 i1_4_lut_adj_45 (.A(n18763), .B(n18756), .C(n18612), .D(n10337), 
         .Z(n34)) /* synthesis lut_function=(A+!(B (C+(D))+!B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(296[16:51])
    defparam i1_4_lut_adj_45.init = 16'habaf;
    LUT4 mux_1597_i1_3_lut (.A(count1[14]), .B(count2[14]), .C(n3064), 
         .Z(n2508[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i1_3_lut.init = 16'hcaca;
    LUT4 i7326_2_lut (.A(count12[14]), .B(n3062), .Z(n2479[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7326_2_lut.init = 16'h8888;
    LUT4 i12200_3_lut (.A(n2595[14]), .B(n2624[14]), .C(n3080), .Z(n2744[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12200_3_lut.init = 16'hcaca;
    PFUMX mux_1604_i6 (.BLUT(n3600[19]), .ALUT(n3573[19]), .C0(n3599), 
          .Z(n3654[19]));
    LUT4 i7615_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[13]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7615_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_2_lut_rep_481_4_lut (.A(n18722), .B(n18813), .C(n6_adj_13), 
         .D(n879), .Z(n18663)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(445[16:65])
    defparam i1_2_lut_rep_481_4_lut.init = 16'hffa2;
    PFUMX mux_1604_i5 (.BLUT(n3600[18]), .ALUT(n3573[18]), .C0(n3599), 
          .Z(n3654[18]));
    LUT4 i7714_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[14]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7714_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1597_i2_3_lut (.A(count1[15]), .B(count2[15]), .C(n3064), 
         .Z(n2508[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i2_3_lut.init = 16'hcaca;
    LUT4 i7551_2_lut (.A(count12[15]), .B(n3062), .Z(n2479[15])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7551_2_lut.init = 16'h8888;
    LUT4 mux_1597_i3_3_lut (.A(count1[16]), .B(count2[16]), .C(n3064), 
         .Z(n2508[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i3_3_lut.init = 16'hcaca;
    LUT4 i7552_2_lut (.A(count12[16]), .B(n3062), .Z(n2479[16])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7552_2_lut.init = 16'h8888;
    PFUMX mux_1604_i4 (.BLUT(n3600[17]), .ALUT(n3573[17]), .C0(n3599), 
          .Z(n3654[17]));
    LUT4 mux_1605_i8_3_lut (.A(count1[21]), .B(count3[21]), .C(\rom2[1] ), 
         .Z(n3371[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1597_i4_3_lut (.A(count1[17]), .B(count2[17]), .C(n3064), 
         .Z(n2508[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i4_3_lut.init = 16'hcaca;
    LUT4 i7553_2_lut (.A(count12[17]), .B(n3062), .Z(n2479[17])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7553_2_lut.init = 16'h8888;
    FD1P3AX en_1__421 (.D(en_1__N_194), .SP(clk_N_168_enable_524), .CK(clk_N_168), 
            .Q(en[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=3, LSE_LLINE=36, LSE_RLINE=45 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(370[8] 432[5])
    defparam en_1__421.GSR = "DISABLED";
    LUT4 mux_1597_i5_3_lut (.A(count1[18]), .B(count2[18]), .C(n3064), 
         .Z(n2508[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i5_3_lut.init = 16'hcaca;
    LUT4 i7554_2_lut (.A(count12[18]), .B(n3062), .Z(n2479[18])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7554_2_lut.init = 16'h8888;
    PFUMX mux_1604_i3 (.BLUT(n3600[16]), .ALUT(n3573[16]), .C0(n3599), 
          .Z(n3654[16]));
    LUT4 mux_1597_i6_3_lut (.A(count1[19]), .B(count2[19]), .C(n3064), 
         .Z(n2508[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i6_3_lut.init = 16'hcaca;
    LUT4 i7555_2_lut (.A(count12[19]), .B(n3062), .Z(n2479[19])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7555_2_lut.init = 16'h8888;
    PFUMX mux_1604_i2 (.BLUT(n3600[15]), .ALUT(n3573[15]), .C0(n3599), 
          .Z(n3654[15]));
    LUT4 mux_1597_i7_3_lut (.A(count1[20]), .B(count2[20]), .C(n3064), 
         .Z(n2508[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i7_3_lut.init = 16'hcaca;
    LUT4 i7556_2_lut (.A(count12[20]), .B(n3062), .Z(n2479[20])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7556_2_lut.init = 16'h8888;
    LUT4 mux_1597_i8_3_lut (.A(count1[21]), .B(count2[21]), .C(n3064), 
         .Z(n2508[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i8_3_lut.init = 16'hcaca;
    LUT4 i7557_2_lut (.A(count12[21]), .B(n3062), .Z(n2479[21])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7557_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_424_3_lut_4_lut_4_lut (.A(n18667), .B(n18685), .C(n18720), 
         .D(n18709), .Z(n18606)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_2_lut_rep_424_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 mux_1597_i9_3_lut (.A(count1[22]), .B(count2[22]), .C(n3064), 
         .Z(n2508[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i9_3_lut.init = 16'hcaca;
    LUT4 i7558_2_lut (.A(count12[22]), .B(n3062), .Z(n2479[22])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7558_2_lut.init = 16'h8888;
    LUT4 mux_1608_i3_3_lut (.A(count11[16]), .B(count7[16]), .C(rom2[2]), 
         .Z(n3458[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1597_i10_3_lut (.A(count1[23]), .B(count2[23]), .C(n3064), 
         .Z(n2508[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i10_3_lut.init = 16'hcaca;
    LUT4 i7616_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[14]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7616_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7559_2_lut (.A(count12[23]), .B(n3062), .Z(n2479[23])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7559_2_lut.init = 16'h8888;
    LUT4 mux_1597_i11_3_lut (.A(count1[24]), .B(count2[24]), .C(n3064), 
         .Z(n2508[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1597_i11_3_lut.init = 16'hcaca;
    LUT4 i7560_2_lut (.A(count12[24]), .B(n3062), .Z(n2479[24])) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i7560_2_lut.init = 16'h8888;
    LUT4 mux_1603_i8_3_lut (.A(count2[21]), .B(count6[21]), .C(rom2[2]), 
         .Z(n3400[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i8_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_461_4_lut (.A(n18721), .B(n5), .C(n6_adj_13), .D(n9292), 
         .Z(n18643)) /* synthesis lut_function=(A (B+(C+(D)))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(439[11:60])
    defparam i1_2_lut_rep_461_4_lut.init = 16'hffa8;
    LUT4 i12214_3_lut (.A(n2595[15]), .B(n2624[15]), .C(n3080), .Z(n2744[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12214_3_lut.init = 16'hcaca;
    LUT4 i12216_3_lut (.A(n2595[16]), .B(n2624[16]), .C(n3080), .Z(n2744[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12216_3_lut.init = 16'hcaca;
    LUT4 mux_1609_i7_3_lut (.A(count4[20]), .B(count5[20]), .C(\rom2[0] ), 
         .Z(n3429[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i7_3_lut.init = 16'hcaca;
    LUT4 i12218_3_lut (.A(n2595[17]), .B(n2624[17]), .C(n3080), .Z(n2744[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12218_3_lut.init = 16'hcaca;
    LUT4 i12220_3_lut (.A(n2595[18]), .B(n2624[18]), .C(n3080), .Z(n2744[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12220_3_lut.init = 16'hcaca;
    LUT4 i12222_3_lut (.A(n2595[19]), .B(n2624[19]), .C(n3080), .Z(n2744[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12222_3_lut.init = 16'hcaca;
    LUT4 i12224_3_lut (.A(n2595[20]), .B(n2624[20]), .C(n3080), .Z(n2744[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12224_3_lut.init = 16'hcaca;
    LUT4 i12226_3_lut (.A(n2595[21]), .B(n2624[21]), .C(n3080), .Z(n2744[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12226_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i3_3_lut (.A(count8[16]), .B(count9[16]), .C(\rom2[0] ), 
         .Z(n3487[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i3_3_lut.init = 16'hcaca;
    LUT4 i12228_3_lut (.A(n2595[22]), .B(n2624[22]), .C(n3080), .Z(n2744[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12228_3_lut.init = 16'hcaca;
    LUT4 i12230_3_lut (.A(n2595[23]), .B(n2624[23]), .C(n3080), .Z(n2744[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12230_3_lut.init = 16'hcaca;
    LUT4 i12232_3_lut (.A(n2595[24]), .B(n2624[24]), .C(n3080), .Z(n2744[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam i12232_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_428_4_lut_4_lut (.A(n18667), .B(n18763), .C(n18668), 
         .D(n18761), .Z(n18610)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i2_3_lut_rep_428_4_lut_4_lut.init = 16'hfffd;
    LUT4 mux_1607_i3_3_lut (.A(n3429[16]), .B(count13[16]), .C(\rom2[3] ), 
         .Z(n3573[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i3_3_lut.init = 16'hcaca;
    LUT4 i7617_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[15]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7617_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1609_i6_3_lut (.A(count4[19]), .B(count5[19]), .C(\rom2[0] ), 
         .Z(n3429[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i6_3_lut.init = 16'hcaca;
    LUT4 i7515_2_lut_rep_478_4_lut (.A(n18761), .B(n18814), .C(n12287), 
         .D(n923), .Z(n18660)) /* synthesis lut_function=(A (B+((D)+!C))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(472[16:68])
    defparam i7515_2_lut_rep_478_4_lut.init = 16'hff8a;
    LUT4 mux_1608_i4_3_lut (.A(count11[17]), .B(count7[17]), .C(rom2[2]), 
         .Z(n3458[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i4_3_lut (.A(count8[17]), .B(count9[17]), .C(\rom2[0] ), 
         .Z(n3487[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i4_3_lut (.A(n3429[17]), .B(count13[17]), .C(\rom2[3] ), 
         .Z(n3573[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i4_3_lut.init = 16'hcaca;
    LUT4 i7514_2_lut_rep_479_4_lut (.A(n18771), .B(n18813), .C(n6), .D(n911), 
         .Z(n18661)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(469[16:68])
    defparam i7514_2_lut_rep_479_4_lut.init = 16'hffa2;
    LUT4 key_flag_11__bdd_2_lut (.A(rom2[2]), .B(\key_flag[9] ), .Z(n18591)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam key_flag_11__bdd_2_lut.init = 16'h1111;
    LUT4 i7618_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[16]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7618_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1608_i5_3_lut (.A(count11[18]), .B(count7[18]), .C(rom2[2]), 
         .Z(n3458[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i5_3_lut (.A(count8[18]), .B(count9[18]), .C(\rom2[0] ), 
         .Z(n3487[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i5_3_lut (.A(n3429[18]), .B(count13[18]), .C(\rom2[3] ), 
         .Z(n3573[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1486_i11_3_lut (.A(n2779[24]), .B(n2809[24]), .C(n3086), 
         .Z(u_count1_24__N_142[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1486_i10_3_lut (.A(n2779[23]), .B(n2809[23]), .C(n3086), 
         .Z(u_count1_24__N_142[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1608_i6_3_lut (.A(count11[19]), .B(count7[19]), .C(rom2[2]), 
         .Z(n3458[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1602_i8_3_lut (.A(count12[21]), .B(count10[21]), .C(\rom2[1] ), 
         .Z(n3516[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i8_3_lut.init = 16'hcaca;
    LUT4 i7265_4_lut (.A(n3815), .B(n444), .C(n11464), .D(n18689), .Z(n3830)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(272[13] 300[21])
    defparam i7265_4_lut.init = 16'h3032;
    LUT4 mux_1602_i11_3_lut (.A(count12[24]), .B(count10[24]), .C(\rom2[1] ), 
         .Z(n3516[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i11_3_lut.init = 16'hcaca;
    LUT4 i7619_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[17]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7619_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7260_4_lut (.A(n480), .B(n468), .C(n18699), .D(n18698), .Z(n3800)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(290[13] 300[21])
    defparam i7260_4_lut.init = 16'h3032;
    LUT4 mux_1602_i10_3_lut (.A(count12[23]), .B(count10[23]), .C(\rom2[1] ), 
         .Z(n3516[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i10_3_lut.init = 16'hcaca;
    LUT4 i7620_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[18]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7620_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1610_i8_3_lut (.A(count8[21]), .B(count9[21]), .C(\rom2[0] ), 
         .Z(n3487[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i8_3_lut.init = 16'hcaca;
    LUT4 i7621_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[19]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7621_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i1_3_lut (.A(count1[14]), .B(count3[14]), .C(\rom2[1] ), 
         .Z(n3371[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i1_3_lut.init = 16'hcaca;
    LUT4 i7720_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[20]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7720_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1603_i1_3_lut (.A(count2[14]), .B(count6[14]), .C(rom2[2]), 
         .Z(n3400[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1602_i1_3_lut (.A(count12[14]), .B(count10[14]), .C(\rom2[1] ), 
         .Z(n3516[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_4_lut (.A(n907), .B(n18661), .C(n903), .D(n18660), 
         .Z(n15938)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(463[13] 479[21])
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    LUT4 i7622_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[20]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7622_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1610_i6_3_lut (.A(count8[19]), .B(count9[19]), .C(\rom2[0] ), 
         .Z(n3487[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i6_3_lut.init = 16'hcaca;
    LUT4 i91_2_lut_rep_540 (.A(\key_value[2] ), .B(\key_flag[2] ), .Z(n18722)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[16:49])
    defparam i91_2_lut_rep_540.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_46 (.A(n18713), .B(n9292), .C(n16929), 
         .D(n18663), .Z(n16930)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(482[8:20])
    defparam i1_2_lut_3_lut_4_lut_adj_46.init = 16'hfffe;
    LUT4 i11953_3_lut (.A(\key_flag[5] ), .B(\key_flag[6] ), .C(rom1[0]), 
         .Z(n17244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11953_3_lut.init = 16'hcaca;
    LUT4 i93_3_lut_rep_494_4_lut (.A(\key_value[2] ), .B(\key_flag[2] ), 
         .C(n18724), .D(n12156), .Z(n18676)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[16:49])
    defparam i93_3_lut_rep_494_4_lut.init = 16'h4044;
    LUT4 i1_2_lut_rep_484_3_lut_4_lut (.A(\key_value[2] ), .B(\key_flag[2] ), 
         .C(n18725), .D(n18736), .Z(n18666)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[16:49])
    defparam i1_2_lut_rep_484_3_lut_4_lut.init = 16'hfff4;
    LUT4 i281_3_lut_rep_530_4_lut (.A(\key_value[2] ), .B(\key_flag[2] ), 
         .C(n6_adj_13), .D(n18813), .Z(n18712)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(266[16:49])
    defparam i281_3_lut_rep_530_4_lut.init = 16'h4044;
    LUT4 i11952_3_lut (.A(\key_flag[3] ), .B(\key_flag[4] ), .C(rom1[0]), 
         .Z(n17243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11952_3_lut.init = 16'hcaca;
    LUT4 i158_3_lut (.A(\key_flag[7] ), .B(\key_flag[8] ), .C(rom1[0]), 
         .Z(n163)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam i158_3_lut.init = 16'h3535;
    LUT4 equal_1580_i6_2_lut_rep_542 (.A(rom2[2]), .B(\rom2[3] ), .Z(n18724)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(260[46:60])
    defparam equal_1580_i6_2_lut_rep_542.init = 16'heeee;
    LUT4 i89_3_lut_4_lut (.A(rom2[2]), .B(\rom2[3] ), .C(n18764), .D(n18725), 
         .Z(n436)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(260[46:60])
    defparam i89_3_lut_4_lut.init = 16'hfe00;
    LUT4 i87_2_lut_rep_543 (.A(\key_value[1] ), .B(\key_flag[1] ), .Z(n18725)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(263[16:49])
    defparam i87_2_lut_rep_543.init = 16'h4444;
    LUT4 i4709_2_lut_rep_502_3_lut_4_lut (.A(\key_value[1] ), .B(\key_flag[1] ), 
         .C(\key_flag[2] ), .D(\key_value[2] ), .Z(n18684)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(263[16:49])
    defparam i4709_2_lut_rep_502_3_lut_4_lut.init = 16'h44f4;
    LUT4 mux_1605_i9_3_lut (.A(count1[22]), .B(count3[22]), .C(\rom2[1] ), 
         .Z(n3371[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1603_i9_3_lut (.A(count2[22]), .B(count6[22]), .C(rom2[2]), 
         .Z(n3400[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1486_i9_3_lut (.A(n2779[22]), .B(n2809[22]), .C(n3086), .Z(u_count1_24__N_142[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_500_3_lut_4_lut (.A(\key_value[1] ), .B(\key_flag[1] ), 
         .C(\key_flag[0] ), .D(\key_value[0] ), .Z(n18682)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(263[16:49])
    defparam i1_2_lut_rep_500_3_lut_4_lut.init = 16'h44f4;
    LUT4 i277_3_lut_4_lut (.A(\key_value[1] ), .B(\key_flag[1] ), .C(n6_adj_13), 
         .D(n5_adj_11), .Z(n879)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(263[16:49])
    defparam i277_3_lut_4_lut.init = 16'h4440;
    LUT4 mux_1486_i8_3_lut (.A(n2779[21]), .B(n2809[21]), .C(n3086), .Z(u_count1_24__N_142[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1486_i7_3_lut (.A(n2779[20]), .B(n2809[20]), .C(n3086), .Z(u_count1_24__N_142[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1486_i6_3_lut (.A(n2779[19]), .B(n2809[19]), .C(n3086), .Z(u_count1_24__N_142[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1486_i5_3_lut (.A(n2779[18]), .B(n2809[18]), .C(n3086), .Z(u_count1_24__N_142[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i5_3_lut.init = 16'hcaca;
    LUT4 i7623_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[21]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7623_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_2_lut_3_lut_4_lut_adj_47 (.A(n9292), .B(n18679), .C(n16816), 
         .D(n18665), .Z(n16916)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(272[13] 300[21])
    defparam i1_2_lut_3_lut_4_lut_adj_47.init = 16'hfffe;
    LUT4 i1_4_lut_adj_48 (.A(n18754), .B(n18667), .C(n18668), .D(n16828), 
         .Z(n358[14])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(290[16:51])
    defparam i1_4_lut_adj_48.init = 16'hc4c0;
    LUT4 i7624_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[22]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7624_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n18667), .B(n18707), .C(n18706), .D(n18668), 
         .Z(n16_adj_1086)) /* synthesis lut_function=((B (D)+!B ((D)+!C))+!A) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hff57;
    LUT4 i11950_3_lut (.A(\key_value[5] ), .B(\key_value[6] ), .C(rom1[0]), 
         .Z(n17241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11950_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_434_4_lut_4_lut (.A(n18667), .B(n16888), .C(n18709), 
         .D(n18668), .Z(n18616)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i2_3_lut_rep_434_4_lut_4_lut.init = 16'hfffd;
    LUT4 mux_1486_i4_3_lut (.A(n2779[17]), .B(n2809[17]), .C(n3086), .Z(u_count1_24__N_142[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i4_3_lut.init = 16'hcaca;
    LUT4 i11949_3_lut (.A(\key_value[3] ), .B(\key_value[4] ), .C(rom1[0]), 
         .Z(n17240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i11949_3_lut.init = 16'hcaca;
    LUT4 i7304_2_lut (.A(\rom2[0] ), .B(\rom2[1] ), .Z(n12156)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7304_2_lut.init = 16'h8888;
    LUT4 i7625_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[23]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7625_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1486_i3_3_lut (.A(n2779[16]), .B(n2809[16]), .C(n3086), .Z(u_count1_24__N_142[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i6_3_lut (.A(n3429[19]), .B(count13[19]), .C(\rom2[3] ), 
         .Z(n3573[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i6_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_550 (.A(\note[1] ), .B(\note[0] ), .Z(n18732)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i2_2_lut_rep_550.init = 16'h2222;
    LUT4 i7626_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[24]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7626_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i4515_4_lut_4_lut_4_lut_4_lut (.A(\note[1] ), .B(\note[0] ), .C(n18807), 
         .D(n18808), .Z(\cycle_17__N_740[3] )) /* synthesis lut_function=(A (B (D)+!B !(C+(D)))+!A (B (D))) */ ;
    defparam i4515_4_lut_4_lut_4_lut_4_lut.init = 16'hcc02;
    LUT4 mux_1486_i2_3_lut (.A(n2779[15]), .B(n2809[15]), .C(n3086), .Z(u_count1_24__N_142[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(313[3] 331[7])
    defparam mux_1486_i2_3_lut.init = 16'hcaca;
    LUT4 i7639_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[13]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7639_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i39_4_lut_then_4_lut (.A(\note[1] ), .B(\note[0] ), .C(n18807), 
         .D(n18808), .Z(n18852)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam i39_4_lut_then_4_lut.init = 16'hf008;
    LUT4 i39_4_lut_else_4_lut (.A(rom1[2]), .B(rom1[3]), .C(rom1[0]), 
         .D(rom1[1]), .Z(n18851)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A !(B))) */ ;
    defparam i39_4_lut_else_4_lut.init = 16'h64c4;
    LUT4 i1_4_lut_adj_49 (.A(n18771), .B(n8), .C(n18720), .D(n18754), 
         .Z(n4)) /* synthesis lut_function=(A+!(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_49.init = 16'hafae;
    PFUMX i12602 (.BLUT(n18817), .ALUT(n18818), .C0(n19846), .Z(n3064));
    LUT4 i7638_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[12]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7638_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_3_lut_rep_555 (.A(\note[3] ), .B(\note[1] ), .C(\note[2] ), 
         .Z(n18737)) /* synthesis lut_function=(A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(335[11:18])
    defparam i1_3_lut_rep_555.init = 16'ha8a8;
    LUT4 i7805_3_lut_4_lut (.A(\note[3] ), .B(\note[1] ), .C(\note[2] ), 
         .D(\note[0] ), .Z(n3_adj_858)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(335[11:18])
    defparam i7805_3_lut_4_lut.init = 16'h3320;
    LUT4 mux_63_Mux_9_i3_3_lut_3_lut_4_lut (.A(\note[3] ), .B(\note[1] ), 
         .C(\note[2] ), .D(\note[0] ), .Z(n3)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (B (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(335[11:18])
    defparam mux_63_Mux_9_i3_3_lut_3_lut_4_lut.init = 16'hcc20;
    LUT4 mux_1608_i7_3_lut (.A(count11[20]), .B(count7[20]), .C(rom2[2]), 
         .Z(n3458[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i7_3_lut.init = 16'hcaca;
    LUT4 i7808_3_lut_4_lut (.A(\note[3] ), .B(\note[1] ), .C(\note[2] ), 
         .D(\note[0] ), .Z(n3_adj_15)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(335[11:18])
    defparam i7808_3_lut_4_lut.init = 16'hff20;
    LUT4 i7802_2_lut_rep_474_3_lut_4_lut (.A(\note[3] ), .B(\note[1] ), 
         .C(\note[2] ), .D(\note[0] ), .Z(n18656)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(335[11:18])
    defparam i7802_2_lut_rep_474_3_lut_4_lut.init = 16'hccec;
    LUT4 i7581_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[4]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7581_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7776_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[14]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7776_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7745_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[20]), .C(\key_value[4] ), 
         .Z(n52[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7745_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7744_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[19]), .C(\key_value[4] ), 
         .Z(n52[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7744_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7775_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[13]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7775_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7743_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[18]), .C(\key_value[4] ), 
         .Z(n52[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7743_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7764_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[2]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[2])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7764_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7742_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[17]), .C(\key_value[4] ), 
         .Z(n52[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7742_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i18_4_lut_4_lut (.A(n19846), .B(n18803), .C(n10301), .D(n18808), 
         .Z(n3066)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(C))) */ ;
    defparam i18_4_lut_4_lut.init = 16'h50d8;
    LUT4 note_4__bdd_4_lut (.A(\note[4] ), .B(\note[3] ), .C(n18803), 
         .D(\note[2] ), .Z(\yinjie_box_2__N_394[0] )) /* synthesis lut_function=(A (B ((D)+!C))+!A ((C+!(D))+!B)) */ ;
    defparam note_4__bdd_4_lut.init = 16'hd95d;
    LUT4 i7741_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[16]), .C(\key_value[4] ), 
         .Z(n52[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7741_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i36_4_lut_4_lut_adj_50 (.A(n19846), .B(n18808), .C(n16871), .D(n18769), 
         .Z(n3078)) /* synthesis lut_function=(!(A (B+!(D))+!A !(C))) */ ;
    defparam i36_4_lut_4_lut_adj_50.init = 16'h7250;
    LUT4 i16_4_lut_4_lut (.A(n19846), .B(n18732), .C(n16843), .D(n18659), 
         .Z(n3072)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;
    defparam i16_4_lut_4_lut.init = 16'hd850;
    LUT4 i7637_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[11]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7637_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7582_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[5]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7582_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i12253_3_lut_4_lut_4_lut (.A(n19846), .B(n414), .C(n18808), .D(n18734), 
         .Z(\cycle_17__N_740[4] )) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam i12253_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i7772_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[10]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7772_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i16_4_lut_4_lut_adj_51 (.A(n19846), .B(n18732), .C(n4_adj_1099), 
         .D(n18808), .Z(n3068)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(C))) */ ;
    defparam i16_4_lut_4_lut_adj_51.init = 16'h50d8;
    LUT4 i1_2_lut (.A(\rom2[0] ), .B(\rom2[1] ), .Z(n5_adj_17)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 mux_63_Mux_16_i15_3_lut_3_lut (.A(n19846), .B(n18610), .C(n18808), 
         .Z(\cycle_17__N_740[16] )) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_63_Mux_16_i15_3_lut_3_lut.init = 16'he4e4;
    LUT4 i12251_3_lut_4_lut_4_lut (.A(n19846), .B(n405), .C(n18732), .D(n18808), 
         .Z(\cycle_17__N_740[13] )) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam i12251_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i7774_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[12]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7774_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7777_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[15]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7777_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1610_i7_3_lut (.A(count8[20]), .B(count9[20]), .C(\rom2[0] ), 
         .Z(n3487[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i7_3_lut.init = 16'hcaca;
    LUT4 i7779_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[17]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7779_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7748_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[23]), .C(\key_value[4] ), 
         .Z(n52[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7748_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7780_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[18]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7780_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1607_i7_3_lut (.A(n3429[20]), .B(count13[20]), .C(\rom2[3] ), 
         .Z(n3573[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i7_3_lut.init = 16'hcaca;
    LUT4 i7778_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[16]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7778_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_63_Mux_9_i15_4_lut_4_lut (.A(n19846), .B(n18610), .C(n262), 
         .D(n18808), .Z(\cycle_17__N_740[9] )) /* synthesis lut_function=(A (D)+!A (B+(C))) */ ;
    defparam mux_63_Mux_9_i15_4_lut_4_lut.init = 16'hfe54;
    LUT4 i7733_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[8]), .C(\key_value[4] ), 
         .Z(n52[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7733_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7726_3_lut_4_lut_4_lut (.A(n19846), .B(count5[1]), .C(fcw_r_adj_1412[0]), 
         .D(\key_value[4] ), .Z(n52[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7726_3_lut_4_lut_4_lut.init = 16'h283c;
    LUT4 i7770_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[8]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7770_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7734_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[9]), .C(\key_value[4] ), 
         .Z(n52[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7734_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7732_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[7]), .C(\key_value[4] ), 
         .Z(n52[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7732_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7721_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[21]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7721_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7715_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[15]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7715_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7728_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[3]), .C(\key_value[4] ), 
         .Z(n52[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7728_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7765_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1404[3]), 
         .C(\key_value[1] ), .Z(n52_adj_1405[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7765_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7730_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[5]), .C(\key_value[4] ), 
         .Z(n52[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7730_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7591_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[14]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7591_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7592_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[15]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7592_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7593_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[16]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7593_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7594_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[17]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7594_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7595_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[18]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7595_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7596_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[19]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7596_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7597_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[20]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7597_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7598_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[21]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7598_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7599_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[22]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7599_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7600_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[23]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7600_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7601_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1406[24]), 
         .C(\key_value[12] ), .Z(n52_adj_1407[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7601_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1609_i5_3_lut (.A(count4[18]), .B(count5[18]), .C(\rom2[0] ), 
         .Z(n3429[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i5_3_lut.init = 16'hcaca;
    LUT4 i7603_3_lut_4_lut_4_lut (.A(n19846), .B(count11[1]), .C(fcw_r_adj_1425[6]), 
         .D(\key_value[10] ), .Z(n52_adj_1401[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7603_3_lut_4_lut_4_lut.init = 16'h283c;
    LUT4 i7604_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[2]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[2])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7604_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7605_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[3]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7605_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7606_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[4]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7606_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7731_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[6]), .C(\key_value[4] ), 
         .Z(n52[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7731_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7727_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[2]), .C(\key_value[4] ), 
         .Z(n52[2])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7727_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7729_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543[4]), .C(\key_value[4] ), 
         .Z(n52[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7729_2_lut_3_lut_3_lut.init = 16'h8c8c;
    CCU2D add_2219_12 (.A0(data_out1[10]), .B0(data_out2[10]), .C0(GND_net), 
          .D0(GND_net), .A1(data_out1[11]), .B1(data_out2[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15481), .COUT(n15482), .S0(\PWM_in_12__N_452[10] ), 
          .S1(\PWM_in_12__N_452[11] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_12.INIT0 = 16'h5666;
    defparam add_2219_12.INIT1 = 16'h5666;
    defparam add_2219_12.INJECT1_0 = "NO";
    defparam add_2219_12.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(rom2[2]), .B(\rom2[3] ), .C(\rom2[1] ), .D(\rom2[0] ), 
         .Z(n3599)) /* synthesis lut_function=(!((B (C+!(D))+!B (C))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(434[1] 485[5])
    defparam i2_4_lut.init = 16'h0a02;
    LUT4 i7608_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[6]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7608_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7636_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[10]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7636_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1609_i8_3_lut (.A(count4[21]), .B(count5[21]), .C(\rom2[0] ), 
         .Z(n3429[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i8_3_lut.init = 16'hcaca;
    CCU2D add_2219_10 (.A0(data_out1[8]), .B0(data_out2[8]), .C0(GND_net), 
          .D0(GND_net), .A1(data_out1[9]), .B1(data_out2[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15480), .COUT(n15481), .S0(\PWM_in_12__N_452[8] ), 
          .S1(\PWM_in_12__N_452[9] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_10.INIT0 = 16'h5666;
    defparam add_2219_10.INIT1 = 16'h5666;
    defparam add_2219_10.INJECT1_0 = "NO";
    defparam add_2219_10.INJECT1_1 = "NO";
    LUT4 i7635_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[9]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7635_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7716_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[16]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7716_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7287_4_lut (.A(n3890[0]), .B(n18677), .C(n903), .D(n907), 
         .Z(n3905[0])) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(460[13] 479[21])
    defparam i7287_4_lut.init = 16'hcfce;
    CCU2D add_2219_8 (.A0(data_out1[6]), .B0(data_out2[6]), .C0(GND_net), 
          .D0(GND_net), .A1(data_out1[7]), .B1(data_out2[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15479), .COUT(n15480), .S0(\PWM_in_12__N_452[6] ), 
          .S1(\PWM_in_12__N_452[7] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_8.INIT0 = 16'h5666;
    defparam add_2219_8.INIT1 = 16'h5666;
    defparam add_2219_8.INJECT1_0 = "NO";
    defparam add_2219_8.INJECT1_1 = "NO";
    LUT4 i7634_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[8]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7634_2_lut_3_lut_3_lut.init = 16'h8c8c;
    CCU2D add_2219_6 (.A0(data_out1[4]), .B0(data_out2[4]), .C0(GND_net), 
          .D0(GND_net), .A1(data_out1[5]), .B1(data_out2[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15478), .COUT(n15479), .S0(\PWM_in_12__N_452[4] ), 
          .S1(\PWM_in_12__N_452[5] ));   // d:/fpga_project/lattice_diamond/piano/speaker.v(554[16:47])
    defparam add_2219_6.INIT0 = 16'h5666;
    defparam add_2219_6.INIT1 = 16'h5666;
    defparam add_2219_6.INJECT1_0 = "NO";
    defparam add_2219_6.INJECT1_1 = "NO";
    LUT4 i7633_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[7]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7633_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7632_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[6]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7632_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7607_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1400[5]), 
         .C(\key_value[10] ), .Z(n52_adj_1401[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7607_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7631_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[5]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7631_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_2_lut_adj_52 (.A(\rom2[1] ), .B(rom2[2]), .Z(n58)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_52.init = 16'h8888;
    LUT4 i7630_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[4]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7630_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7629_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[3]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7629_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7628_3_lut_4_lut_4_lut (.A(n19846), .B(count10[2]), .C(fcw_r_adj_1426[2]), 
         .D(\key_value[9] ), .Z(n52_adj_1424[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7628_3_lut_4_lut_4_lut.init = 16'h283c;
    LUT4 i7640_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[14]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7640_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7641_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[15]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7641_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7642_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[16]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7642_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7643_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[17]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7643_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7644_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[18]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7644_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1609_i4_3_lut (.A(count4[17]), .B(count5[17]), .C(\rom2[0] ), 
         .Z(n3429[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i4_3_lut.init = 16'hcaca;
    LUT4 i7283_4_lut (.A(n923), .B(n911), .C(n18719), .D(n18718), .Z(n3890[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(469[13] 479[21])
    defparam i7283_4_lut.init = 16'h3032;
    LUT4 i7645_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[19]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7645_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7646_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[20]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7646_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7647_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[21]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7647_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7648_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[22]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7648_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7649_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[23]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7649_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7650_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1423[24]), 
         .C(\key_value[9] ), .Z(n52_adj_1424[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7650_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7652_3_lut_4_lut_4_lut (.A(n19846), .B(count9[1]), .C(fcw_r_adj_1427[8]), 
         .D(\key_value[8] ), .Z(n52_adj_1428[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7652_3_lut_4_lut_4_lut.init = 16'h283c;
    LUT4 key_flag_11__bdd_3_lut (.A(\key_flag[11] ), .B(rom2[2]), .C(\key_flag[7] ), 
         .Z(n18592)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+!(C)))) */ ;
    defparam key_flag_11__bdd_3_lut.init = 16'h4747;
    LUT4 i7653_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[2]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[2])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7653_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7654_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[3]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7654_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7655_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[4]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7655_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7656_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[5]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7656_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7657_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[6]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7657_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7658_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[7]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7658_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7659_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[8]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7659_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7660_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[9]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7660_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7661_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[10]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7661_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7662_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[11]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7662_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_4_lut_adj_53 (.A(n18768), .B(n18685), .C(n18720), .D(n31), 
         .Z(n351)) /* synthesis lut_function=(!(A+!(B+!(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(287[16:49])
    defparam i1_4_lut_adj_53.init = 16'h4544;
    LUT4 i7663_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[12]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7663_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7664_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[13]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7664_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7665_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[14]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7665_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7666_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[15]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7666_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7667_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[16]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7667_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7668_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[17]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7668_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX mux_1604_i1 (.BLUT(n3600[14]), .ALUT(n3573[14]), .C0(n3599), 
          .Z(n3654[14]));
    LUT4 i7669_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[18]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7669_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7670_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[19]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7670_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7671_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[20]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7671_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7672_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[21]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7672_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7673_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[22]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7673_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1608_i9_3_lut (.A(count11[22]), .B(count7[22]), .C(rom2[2]), 
         .Z(n3458[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i9_3_lut.init = 16'hcaca;
    LUT4 i7674_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[23]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7674_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7675_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1429[24]), 
         .C(\key_value[8] ), .Z(n52_adj_1428[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7675_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1602_i9_3_lut (.A(count12[22]), .B(count10[22]), .C(\rom2[1] ), 
         .Z(n3516[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i9_3_lut.init = 16'hcaca;
    PFUMX i12626 (.BLUT(n18854), .ALUT(n18855), .C0(rom2[2]), .Z(n18856));
    LUT4 mux_1610_i9_3_lut (.A(count8[22]), .B(count9[22]), .C(\rom2[0] ), 
         .Z(n3487[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1264_i1_3_lut (.A(\key_value[11] ), .B(\key_value[12] ), .C(rom1[0]), 
         .Z(n10879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(194[3] 249[17])
    defparam mux_1264_i1_3_lut.init = 16'hcaca;
    LUT4 i7688_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[12]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[12])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7688_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i3_4_lut_adj_54 (.A(n18666), .B(n18655), .C(n18680), .D(n18611), 
         .Z(clk_N_168_enable_507)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[16:49])
    defparam i3_4_lut_adj_54.init = 16'hfffe;
    LUT4 mux_1607_i9_3_lut (.A(n3429[22]), .B(count13[22]), .C(\rom2[3] ), 
         .Z(n3573[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1608_i10_3_lut (.A(count11[23]), .B(count7[23]), .C(rom2[2]), 
         .Z(n3458[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i10_3_lut (.A(count8[23]), .B(count9[23]), .C(\rom2[0] ), 
         .Z(n3487[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i10_3_lut.init = 16'hcaca;
    LUT4 i7687_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[11]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[11])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7687_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7717_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[17]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7717_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1607_i10_3_lut (.A(n3429[23]), .B(count13[23]), .C(\rom2[3] ), 
         .Z(n3573[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i10_3_lut.init = 16'hcaca;
    LUT4 i7686_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[10]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[10])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7686_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1608_i11_3_lut (.A(count11[24]), .B(count7[24]), .C(rom2[2]), 
         .Z(n3458[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1608_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1610_i11_3_lut (.A(count8[24]), .B(count9[24]), .C(\rom2[0] ), 
         .Z(n3487[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1610_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1607_i11_3_lut (.A(n3429[24]), .B(count13[24]), .C(\rom2[3] ), 
         .Z(n3573[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1607_i11_3_lut.init = 16'hcaca;
    LUT4 i7722_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[22]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7722_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7685_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[9]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7685_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7684_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[8]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7684_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7683_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[7]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7683_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7682_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[6]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7682_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 n16967_bdd_3_lut_then_3_lut (.A(\key_flag[4] ), .B(\key_flag[12] ), 
         .C(\rom2[3] ), .Z(n18855)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n16967_bdd_3_lut_then_3_lut.init = 16'h3535;
    LUT4 i7681_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[5]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7681_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1609_i3_3_lut (.A(count4[16]), .B(count5[16]), .C(\rom2[0] ), 
         .Z(n3429[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1609_i3_3_lut.init = 16'hcaca;
    LUT4 i7680_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[4]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7680_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7679_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[3]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7679_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i2_3_lut (.A(count1[15]), .B(count3[15]), .C(\rom2[1] ), 
         .Z(n3371[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i2_3_lut.init = 16'hcaca;
    LUT4 i7678_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[2]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[2])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7678_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX mux_1600_i2 (.BLUT(n3546[15]), .ALUT(n3516[15]), .C0(\rom2[3] ), 
          .Z(n3627[15]));
    LUT4 i7677_3_lut_4_lut_4_lut (.A(n19846), .B(count8[1]), .C(fcw_r_adj_1432[8]), 
         .D(\key_value[7] ), .Z(n52_adj_1431[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7677_3_lut_4_lut_4_lut.init = 16'h283c;
    LUT4 mux_1603_i2_3_lut (.A(count2[15]), .B(count6[15]), .C(rom2[2]), 
         .Z(n3400[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1602_i2_3_lut (.A(count12[15]), .B(count10[15]), .C(\rom2[1] ), 
         .Z(n3516[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i2_3_lut.init = 16'hcaca;
    LUT4 i7689_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[13]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[13])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7689_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i3_3_lut (.A(count1[16]), .B(count3[16]), .C(\rom2[1] ), 
         .Z(n3371[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i3_3_lut.init = 16'hcaca;
    PFUMX mux_1600_i3 (.BLUT(n3546[16]), .ALUT(n3516[16]), .C0(\rom2[3] ), 
          .Z(n3627[16]));
    LUT4 i7690_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[14]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[14])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7690_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7691_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[15]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[15])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7691_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX i11951 (.BLUT(n17240), .ALUT(n17241), .C0(rom1[1]), .Z(n17242));
    PFUMX mux_1600_i4 (.BLUT(n3546[17]), .ALUT(n3516[17]), .C0(\rom2[3] ), 
          .Z(n3627[17]));
    LUT4 mux_1603_i3_3_lut (.A(count2[16]), .B(count6[16]), .C(rom2[2]), 
         .Z(n3400[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i3_3_lut.init = 16'hcaca;
    LUT4 i7692_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[16]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[16])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7692_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX mux_1600_i5 (.BLUT(n3546[18]), .ALUT(n3516[18]), .C0(\rom2[3] ), 
          .Z(n3627[18]));
    LUT4 mux_1602_i3_3_lut (.A(count12[16]), .B(count10[16]), .C(\rom2[1] ), 
         .Z(n3516[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i3_3_lut.init = 16'hcaca;
    PFUMX mux_1600_i6 (.BLUT(n3546[19]), .ALUT(n3516[19]), .C0(\rom2[3] ), 
          .Z(n3627[19]));
    LUT4 i7693_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[17]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[17])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7693_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7694_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[18]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[18])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7694_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i4_3_lut (.A(count1[17]), .B(count3[17]), .C(\rom2[1] ), 
         .Z(n3371[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i4_3_lut.init = 16'hcaca;
    PFUMX mux_1600_i7 (.BLUT(n3546[20]), .ALUT(n3516[20]), .C0(\rom2[3] ), 
          .Z(n3627[20]));
    LUT4 i7695_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[19]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[19])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7695_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1603_i4_3_lut (.A(count2[17]), .B(count6[17]), .C(rom2[2]), 
         .Z(n3400[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i4_3_lut.init = 16'hcaca;
    LUT4 i7696_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[20]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[20])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7696_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7697_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[21]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[21])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7697_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1602_i4_3_lut (.A(count12[17]), .B(count10[17]), .C(\rom2[1] ), 
         .Z(n3516[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i4_3_lut.init = 16'hcaca;
    PFUMX mux_1600_i8 (.BLUT(n3546[21]), .ALUT(n3516[21]), .C0(\rom2[3] ), 
          .Z(n3627[21]));
    LUT4 mux_1605_i5_3_lut (.A(count1[18]), .B(count3[18]), .C(\rom2[1] ), 
         .Z(n3371[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1603_i5_3_lut (.A(count2[18]), .B(count6[18]), .C(rom2[2]), 
         .Z(n3400[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i5_3_lut.init = 16'hcaca;
    LUT4 i7698_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[22]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[22])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7698_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX mux_1600_i9 (.BLUT(n3546[22]), .ALUT(n3516[22]), .C0(\rom2[3] ), 
          .Z(n3627[22]));
    LUT4 i7699_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[23]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[23])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7699_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7700_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1430[24]), 
         .C(\key_value[7] ), .Z(n52_adj_1431[24])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7700_2_lut_3_lut_3_lut.init = 16'h8c8c;
    PFUMX mux_1600_i10 (.BLUT(n3546[23]), .ALUT(n3516[23]), .C0(\rom2[3] ), 
          .Z(n3627[23]));
    LUT4 mux_1602_i5_3_lut (.A(count12[18]), .B(count10[18]), .C(\rom2[1] ), 
         .Z(n3516[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i5_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_55 (.A(n18653), .B(n16876), .C(n18720), .D(n16917), 
         .Z(clk_N_168_enable_518)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(269[16:49])
    defparam i3_4_lut_adj_55.init = 16'hfffe;
    LUT4 i7702_3_lut_4_lut_4_lut (.A(n19846), .B(count6[2]), .C(fcw_r_adj_1412[0]), 
         .D(\key_value[5] ), .Z(n52_adj_1403[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+(D))+!B ((D)+!C)))) */ ;
    defparam i7702_3_lut_4_lut_4_lut.init = 16'h283c;
    PFUMX mux_1600_i11 (.BLUT(n3546[24]), .ALUT(n3516[24]), .C0(\rom2[3] ), 
          .Z(n3627[24]));
    LUT4 i7703_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[3]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7703_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7704_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[4]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[4])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7704_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7705_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[5]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[5])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7705_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1605_i6_3_lut (.A(count1[19]), .B(count3[19]), .C(\rom2[1] ), 
         .Z(n3371[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i6_3_lut.init = 16'hcaca;
    LUT4 i7706_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[6]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[6])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7706_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1603_i6_3_lut (.A(count2[19]), .B(count6[19]), .C(rom2[2]), 
         .Z(n3400[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1603_i6_3_lut.init = 16'hcaca;
    LUT4 i7707_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[7]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[7])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7707_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7708_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[8]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[8])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7708_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 i7709_2_lut_3_lut_3_lut (.A(n19846), .B(count_24__N_543_adj_1402[9]), 
         .C(\key_value[5] ), .Z(n52_adj_1403[9])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i7709_2_lut_3_lut_3_lut.init = 16'h8c8c;
    LUT4 mux_1602_i6_3_lut (.A(count12[19]), .B(count10[19]), .C(\rom2[1] ), 
         .Z(n3516[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1602_i6_3_lut.init = 16'hcaca;
    PFUMX i11945 (.BLUT(n17234), .ALUT(n17235), .C0(\rom2[1] ), .Z(n17236));
    PFUMX mux_1600_i1 (.BLUT(n3546[14]), .ALUT(n3516[14]), .C0(\rom2[3] ), 
          .Z(n3627[14]));
    LUT4 mux_1605_i10_3_lut (.A(count1[23]), .B(count3[23]), .C(\rom2[1] ), 
         .Z(n3371[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_1605_i10_3_lut.init = 16'hcaca;
    DDS u_DDS_9 (.\fcw_r[8] (fcw_r_adj_1427[8]), .clk_N_168(clk_N_168), 
        .n18785(n18785), .\count9[23] (count9[23]), .GND_net(GND_net), 
        .\count9[24] (count9[24]), .\count_24__N_543[23] (count_24__N_543_adj_1429[23]), 
        .\count_24__N_543[24] (count_24__N_543_adj_1429[24]), .\count9[21] (count9[21]), 
        .\count9[22] (count9[22]), .\count_24__N_543[21] (count_24__N_543_adj_1429[21]), 
        .\count_24__N_543[22] (count_24__N_543_adj_1429[22]), .\count9[19] (count9[19]), 
        .\count9[20] (count9[20]), .\count_24__N_543[19] (count_24__N_543_adj_1429[19]), 
        .\count_24__N_543[20] (count_24__N_543_adj_1429[20]), .\count9[17] (count9[17]), 
        .\count9[18] (count9[18]), .\count_24__N_543[17] (count_24__N_543_adj_1429[17]), 
        .\count_24__N_543[18] (count_24__N_543_adj_1429[18]), .\count9[15] (count9[15]), 
        .\count9[16] (count9[16]), .\count_24__N_543[15] (count_24__N_543_adj_1429[15]), 
        .\count_24__N_543[16] (count_24__N_543_adj_1429[16]), .\count9[14] (count9[14]), 
        .\count_24__N_543[13] (count_24__N_543_adj_1429[13]), .\count_24__N_543[14] (count_24__N_543_adj_1429[14]), 
        .\count_24__N_543[11] (count_24__N_543_adj_1429[11]), .\count_24__N_543[12] (count_24__N_543_adj_1429[12]), 
        .\count_24__N_543[9] (count_24__N_543_adj_1429[9]), .\count_24__N_543[10] (count_24__N_543_adj_1429[10]), 
        .\count_24__N_543[7] (count_24__N_543_adj_1429[7]), .\count_24__N_543[8] (count_24__N_543_adj_1429[8]), 
        .\count_24__N_543[5] (count_24__N_543_adj_1429[5]), .\count_24__N_543[6] (count_24__N_543_adj_1429[6]), 
        .\count_24__N_543[3] (count_24__N_543_adj_1429[3]), .\count_24__N_543[4] (count_24__N_543_adj_1429[4]), 
        .\count9[1] (count9[1]), .\count_24__N_543[2] (count_24__N_543_adj_1429[2]), 
        .pwm_out2_N_125(pwm_out2_N_125), .n49(n52_adj_1428[1]), .n48(n52_adj_1428[2]), 
        .n47(n52_adj_1428[3]), .n46(n52_adj_1428[4]), .n45(n52_adj_1428[5]), 
        .n44(n52_adj_1428[6]), .n43(n52_adj_1428[7]), .n42(n52_adj_1428[8]), 
        .n41(n52_adj_1428[9]), .n40(n52_adj_1428[10]), .n39(n52_adj_1428[11]), 
        .n38(n52_adj_1428[12]), .n37(n52_adj_1428[13]), .n36(n52_adj_1428[14]), 
        .n35(n52_adj_1428[15]), .n34(n52_adj_1428[16]), .n33(n52_adj_1428[17]), 
        .n32(n52_adj_1428[18]), .n31(n52_adj_1428[19]), .n30(n52_adj_1428[20]), 
        .n29(n52_adj_1428[21]), .n28(n52_adj_1428[22]), .n27(n52_adj_1428[23]), 
        .n26(n52_adj_1428[24]), .n18784(n18784), .n18757(n18757)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(135[5] 144[3])
    DDS_U0 u_DDS_8 (.\fcw_r[8] (fcw_r_adj_1432[8]), .clk_N_168(clk_N_168), 
           .n18785(n18785), .\count8[23] (count8[23]), .GND_net(GND_net), 
           .\count8[24] (count8[24]), .\count_24__N_543[23] (count_24__N_543_adj_1430[23]), 
           .\count_24__N_543[24] (count_24__N_543_adj_1430[24]), .\count8[21] (count8[21]), 
           .\count8[22] (count8[22]), .\count_24__N_543[21] (count_24__N_543_adj_1430[21]), 
           .\count_24__N_543[22] (count_24__N_543_adj_1430[22]), .\count8[19] (count8[19]), 
           .\count8[20] (count8[20]), .\count_24__N_543[19] (count_24__N_543_adj_1430[19]), 
           .\count_24__N_543[20] (count_24__N_543_adj_1430[20]), .\count8[17] (count8[17]), 
           .\count8[18] (count8[18]), .\count_24__N_543[17] (count_24__N_543_adj_1430[17]), 
           .\count_24__N_543[18] (count_24__N_543_adj_1430[18]), .\count8[15] (count8[15]), 
           .\count8[16] (count8[16]), .\count_24__N_543[15] (count_24__N_543_adj_1430[15]), 
           .\count_24__N_543[16] (count_24__N_543_adj_1430[16]), .\count8[14] (count8[14]), 
           .\count_24__N_543[13] (count_24__N_543_adj_1430[13]), .\count_24__N_543[14] (count_24__N_543_adj_1430[14]), 
           .\count_24__N_543[11] (count_24__N_543_adj_1430[11]), .\count_24__N_543[12] (count_24__N_543_adj_1430[12]), 
           .\count_24__N_543[9] (count_24__N_543_adj_1430[9]), .\count_24__N_543[10] (count_24__N_543_adj_1430[10]), 
           .\count_24__N_543[7] (count_24__N_543_adj_1430[7]), .\count_24__N_543[8] (count_24__N_543_adj_1430[8]), 
           .\count_24__N_543[5] (count_24__N_543_adj_1430[5]), .\count_24__N_543[6] (count_24__N_543_adj_1430[6]), 
           .\count_24__N_543[3] (count_24__N_543_adj_1430[3]), .\count_24__N_543[4] (count_24__N_543_adj_1430[4]), 
           .\count8[1] (count8[1]), .\count_24__N_543[2] (count_24__N_543_adj_1430[2]), 
           .pwm_out2_N_125(pwm_out2_N_125), .n49(n52_adj_1431[1]), .n48(n52_adj_1431[2]), 
           .n47(n52_adj_1431[3]), .n46(n52_adj_1431[4]), .n45(n52_adj_1431[5]), 
           .n44(n52_adj_1431[6]), .n43(n52_adj_1431[7]), .n42(n52_adj_1431[8]), 
           .n41(n52_adj_1431[9]), .n40(n52_adj_1431[10]), .n39(n52_adj_1431[11]), 
           .n38(n52_adj_1431[12]), .n37(n52_adj_1431[13]), .n36(n52_adj_1431[14]), 
           .n35(n52_adj_1431[15]), .n34(n52_adj_1431[16]), .n33(n52_adj_1431[17]), 
           .n32(n52_adj_1431[18]), .n31(n52_adj_1431[19]), .n30(n52_adj_1431[20]), 
           .n29(n52_adj_1431[21]), .n28(n52_adj_1431[22]), .n27(n52_adj_1431[23]), 
           .n26(n52_adj_1431[24]), .n18784(n18784), .n18757(n18757)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(124[5] 133[3])
    DDS_U1 u_DDS_7 (.clk_N_168(clk_N_168), .n18705(n18705), .\count7[24] (count7[24]), 
           .GND_net(GND_net), .n106(n105_adj_1419[24]), .\count7[22] (count7[22]), 
           .\count7[23] (count7[23]), .n108(n105_adj_1419[22]), .n107(n105_adj_1419[23]), 
           .\count7[20] (count7[20]), .\count7[21] (count7[21]), .n110(n105_adj_1419[20]), 
           .n109(n105_adj_1419[21]), .\count7[18] (count7[18]), .\count7[19] (count7[19]), 
           .n112(n105_adj_1419[18]), .n111(n105_adj_1419[19]), .\count7[16] (count7[16]), 
           .\count7[17] (count7[17]), .n114(n105_adj_1419[16]), .n113(n105_adj_1419[17]), 
           .\count7[14] (count7[14]), .\count7[15] (count7[15]), .n116(n105_adj_1419[14]), 
           .n115(n105_adj_1419[15]), .n118(n105_adj_1419[12]), .n117(n105_adj_1419[13]), 
           .n120(n105_adj_1419[10]), .n119(n105_adj_1419[11]), .\fcw_r[8] (fcw_r_adj_1417[8]), 
           .n122(n105_adj_1419[8]), .n121(n105_adj_1419[9]), .n124(n105_adj_1419[6]), 
           .n123(n105_adj_1419[7]), .n126(n105_adj_1419[4]), .n125(n105_adj_1419[5]), 
           .n128(n105_adj_1419[2]), .n127(n105_adj_1419[3]), .n25(n184_adj_1416[0]), 
           .n129(n105_adj_1419[1]), .pwm_out2_N_125(pwm_out2_N_125), .n132({n132_adj_1418}), 
           .n18717(n18717), .n19839(n19839), .n19840(n19840), .n18785(n18785), 
           .n18784(n18784), .n18757(n18757)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(113[5] 122[3])
    DDS_U2 u_DDS_6 (.\count6[24] (count6[24]), .GND_net(GND_net), .\count_24__N_543[24] (count_24__N_543_adj_1402[24]), 
           .\count6[22] (count6[22]), .\count6[23] (count6[23]), .\count_24__N_543[22] (count_24__N_543_adj_1402[22]), 
           .\count_24__N_543[23] (count_24__N_543_adj_1402[23]), .\count6[20] (count6[20]), 
           .\count6[21] (count6[21]), .\count_24__N_543[20] (count_24__N_543_adj_1402[20]), 
           .\count_24__N_543[21] (count_24__N_543_adj_1402[21]), .\count6[18] (count6[18]), 
           .\count6[19] (count6[19]), .\count_24__N_543[18] (count_24__N_543_adj_1402[18]), 
           .\count_24__N_543[19] (count_24__N_543_adj_1402[19]), .\count6[16] (count6[16]), 
           .\count6[17] (count6[17]), .\count_24__N_543[16] (count_24__N_543_adj_1402[16]), 
           .\count_24__N_543[17] (count_24__N_543_adj_1402[17]), .\count6[14] (count6[14]), 
           .\count6[15] (count6[15]), .\count_24__N_543[14] (count_24__N_543_adj_1402[14]), 
           .\count_24__N_543[15] (count_24__N_543_adj_1402[15]), .\count_24__N_543[12] (count_24__N_543_adj_1402[12]), 
           .\count_24__N_543[13] (count_24__N_543_adj_1402[13]), .\fcw_r[2] (fcw_r_adj_1433[2]), 
           .\count_24__N_543[10] (count_24__N_543_adj_1402[10]), .\count_24__N_543[11] (count_24__N_543_adj_1402[11]), 
           .\fcw_r[1] (fcw_r_adj_1433[1]), .\count_24__N_543[8] (count_24__N_543_adj_1402[8]), 
           .\count_24__N_543[9] (count_24__N_543_adj_1402[9]), .\fcw_r[0] (fcw_r_adj_1412[0]), 
           .\count_24__N_543[6] (count_24__N_543_adj_1402[6]), .\count_24__N_543[7] (count_24__N_543_adj_1402[7]), 
           .\fcw_r[4] (fcw_r_adj_1434[4]), .\count_24__N_543[4] (count_24__N_543_adj_1402[4]), 
           .\count_24__N_543[5] (count_24__N_543_adj_1402[5]), .\count6[2] (count6[2]), 
           .\count_24__N_543[3] (count_24__N_543_adj_1402[3]), .n18717(n18717), 
           .n18634(n18634), .\fcw_r_15__N_495[11] (\fcw_r_15__N_495[11] ), 
           .n19839(n19839), .clk_N_168(clk_N_168), .pwm_out2_N_125(pwm_out2_N_125), 
           .n48(n52_adj_1403[2]), .n47(n52_adj_1403[3]), .n46(n52_adj_1403[4]), 
           .n45(n52_adj_1403[5]), .n44(n52_adj_1403[6]), .n43(n52_adj_1403[7]), 
           .n42(n52_adj_1403[8]), .n41(n52_adj_1403[9]), .n40(n52_adj_1403[10]), 
           .n39(n52_adj_1403[11]), .n38(n52_adj_1403[12]), .n37(n52_adj_1403[13]), 
           .n36(n52_adj_1403[14]), .n35(n52_adj_1403[15]), .n34(n52_adj_1403[16]), 
           .n33(n52_adj_1403[17]), .n32(n52_adj_1403[18]), .n31(n52_adj_1403[19]), 
           .n30(n52_adj_1403[20]), .n29(n52_adj_1403[21]), .n28(n52_adj_1403[22]), 
           .n27(n52_adj_1403[23]), .n26(n52_adj_1403[24]), .\fcw_r_15__N_495[8] (fcw_r_15__N_495[8]), 
           .\fcw_r_15__N_495[5] (\fcw_r_15__N_495[5] ), .n16936(n16936), 
           .n15966(n15966), .n7920(n7919[7])) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(102[5] 111[3])
    DDS_U3 u_DDS_5 (.\count5[23] (count5[23]), .GND_net(GND_net), .\count5[24] (count5[24]), 
           .\count_24__N_543[23] (count_24__N_543[23]), .\count_24__N_543[24] (count_24__N_543[24]), 
           .\count5[21] (count5[21]), .\count5[22] (count5[22]), .\count_24__N_543[21] (count_24__N_543[21]), 
           .\count_24__N_543[22] (count_24__N_543[22]), .\count5[19] (count5[19]), 
           .\count5[20] (count5[20]), .\count_24__N_543[19] (count_24__N_543[19]), 
           .\count_24__N_543[20] (count_24__N_543[20]), .\count5[17] (count5[17]), 
           .\count5[18] (count5[18]), .\count_24__N_543[17] (count_24__N_543[17]), 
           .\count_24__N_543[18] (count_24__N_543[18]), .\count5[15] (count5[15]), 
           .\count5[16] (count5[16]), .\count_24__N_543[15] (count_24__N_543[15]), 
           .\count_24__N_543[16] (count_24__N_543[16]), .\count5[14] (count5[14]), 
           .\count_24__N_543[13] (count_24__N_543[13]), .\count_24__N_543[14] (count_24__N_543[14]), 
           .\fcw_r[1] (fcw_r_adj_1433[1]), .\count_24__N_543[11] (count_24__N_543[11]), 
           .\count_24__N_543[12] (count_24__N_543[12]), .\count5[1] (count5[1]), 
           .clk_N_168(clk_N_168), .pwm_out2_N_125(pwm_out2_N_125), .n49(n52[1]), 
           .n48(n52[2]), .n47(n52[3]), .n46(n52[4]), .n45(n52[5]), .n44(n52[6]), 
           .n43(n52[7]), .n42(n52[8]), .n41(n52[9]), .n40(n52[10]), 
           .n39(n52[11]), .n38(n52[12]), .n37(n52[13]), .n36(n52[14]), 
           .n35(n52[15]), .n34(n52[16]), .n33(n52[17]), .n32(n52[18]), 
           .n31(n52[19]), .n30(n52[20]), .n29(n52[21]), .n28(n52[22]), 
           .n27(n52[23]), .n26(n52[24]), .\fcw_r[2] (fcw_r_adj_1433[2]), 
           .\count_24__N_543[9] (count_24__N_543[9]), .\count_24__N_543[10] (count_24__N_543[10]), 
           .\fcw_r[0] (fcw_r_adj_1412[0]), .\count_24__N_543[7] (count_24__N_543[7]), 
           .\count_24__N_543[8] (count_24__N_543[8]), .n18705(n18705), .n18717(n18717), 
           .n19839(n19839), .n8147(n8147), .n8146(n8146), .n19840(n19840), 
           .\count_24__N_543[5] (count_24__N_543[5]), .\count_24__N_543[6] (count_24__N_543[6]), 
           .\count_24__N_543[3] (count_24__N_543[3]), .\count_24__N_543[4] (count_24__N_543[4]), 
           .\count_24__N_543[2] (count_24__N_543[2])) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(91[5] 100[3])
    DDS_U4 u_DDS_4 (.\fcw_r[1] (fcw_r_adj_1433[1]), .clk_N_168(clk_N_168), 
           .n18784(n18784), .\count4[24] (count4[24]), .GND_net(GND_net), 
           .n106(n105_adj_1413[24]), .\count4[22] (count4[22]), .\count4[23] (count4[23]), 
           .n108(n105_adj_1413[22]), .n107(n105_adj_1413[23]), .\count4[20] (count4[20]), 
           .\count4[21] (count4[21]), .n110(n105_adj_1413[20]), .n109(n105_adj_1413[21]), 
           .\count4[18] (count4[18]), .\count4[19] (count4[19]), .n112(n105_adj_1413[18]), 
           .n111(n105_adj_1413[19]), .\count4[16] (count4[16]), .\count4[17] (count4[17]), 
           .n114(n105_adj_1413[16]), .n113(n105_adj_1413[17]), .\count4[14] (count4[14]), 
           .\count4[15] (count4[15]), .n116(n105_adj_1413[14]), .n115(n105_adj_1413[15]), 
           .n118(n105_adj_1413[12]), .n117(n105_adj_1413[13]), .n120(n105_adj_1413[10]), 
           .n119(n105_adj_1413[11]), .\fcw_r[2] (fcw_r_adj_1433[2]), .n122(n105_adj_1413[8]), 
           .n121(n105_adj_1413[9]), .\fcw_r[0] (fcw_r_adj_1412[0]), .n124(n105_adj_1413[6]), 
           .n123(n105_adj_1413[7]), .n126(n105_adj_1413[4]), .n125(n105_adj_1413[5]), 
           .n128(n105_adj_1413[2]), .n127(n105_adj_1413[3]), .n25(n184_adj_1415[0]), 
           .n129(n105_adj_1413[1]), .pwm_out2_N_125(pwm_out2_N_125), .n132({n132_adj_1414}), 
           .n18757(n18757), .\fcw_r_15__N_495[11] (\fcw_r_15__N_495[11] ), 
           .yinjie({yinjie}), .n18785(n18785), .n19846(n19846), .\yinjie_box[1] (yinjie_box[1]), 
           .\fcw_r_15__N_527[0] (fcw_r_15__N_527[0]), .clk__inv(clk__inv)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(80[5] 89[3])
    DDS_U5 u_DDS_3 (.\fcw_r[0] (fcw_r_adj_1412[0]), .clk_N_168(clk_N_168), 
           .n18785(n18785), .\count3[24] (count3[24]), .GND_net(GND_net), 
           .n106(n105_adj_1409[24]), .\count3[22] (count3[22]), .\count3[23] (count3[23]), 
           .n108(n105_adj_1409[22]), .n107(n105_adj_1409[23]), .\count3[20] (count3[20]), 
           .\count3[21] (count3[21]), .n110(n105_adj_1409[20]), .n109(n105_adj_1409[21]), 
           .\count3[18] (count3[18]), .\count3[19] (count3[19]), .n112(n105_adj_1409[18]), 
           .n111(n105_adj_1409[19]), .\count3[16] (count3[16]), .\count3[17] (count3[17]), 
           .n114(n105_adj_1409[16]), .n113(n105_adj_1409[17]), .\count3[14] (count3[14]), 
           .\count3[15] (count3[15]), .n116(n105_adj_1409[14]), .n115(n105_adj_1409[15]), 
           .n118(n105_adj_1409[12]), .n117(n105_adj_1409[13]), .\fcw_r[2] (fcw_r_adj_1433[2]), 
           .n120(n105_adj_1409[10]), .n119(n105_adj_1409[11]), .\fcw_r[1] (fcw_r_adj_1433[1]), 
           .n122(n105_adj_1409[8]), .n121(n105_adj_1409[9]), .n124(n105_adj_1409[6]), 
           .n123(n105_adj_1409[7]), .n126(n105_adj_1409[4]), .n125(n105_adj_1409[5]), 
           .\fcw_r[4] (fcw_r_adj_1434[4]), .n128(n105_adj_1409[2]), .n127(n105_adj_1409[3]), 
           .n25(n184_adj_1411[0]), .n129(n105_adj_1409[1]), .pwm_out2_N_125(pwm_out2_N_125), 
           .n132({n132_adj_1410}), .\yinjie[2] (yinjie[2]), .n19846(n19846), 
           .n18784(n18784), .\fcw_r_15__N_495[11] (\fcw_r_15__N_495[11] ), 
           .\fcw_r_15__N_495[9] (\fcw_r_15__N_495[9] ), .\fcw_r_15__N_527[0] (fcw_r_15__N_527[0]), 
           .\yinjie[0] (yinjie[0]), .clk__inv(clk__inv)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(69[5] 78[3])
    DDS_U6 u_DDS_2 (.clk_N_168(clk_N_168), .n18784(n18784), .\count2[23] (count2[23]), 
           .GND_net(GND_net), .\count2[24] (count2[24]), .\count_24__N_543[23] (count_24__N_543_adj_1404[23]), 
           .\count_24__N_543[24] (count_24__N_543_adj_1404[24]), .\yinjie[1] (yinjie[1]), 
           .n19846(n19846), .\yinjie[2] (yinjie[2]), .n19840(n19840), 
           .\count2[21] (count2[21]), .\count2[22] (count2[22]), .\count_24__N_543[21] (count_24__N_543_adj_1404[21]), 
           .\count_24__N_543[22] (count_24__N_543_adj_1404[22]), .\count2[19] (count2[19]), 
           .\count2[20] (count2[20]), .\count_24__N_543[19] (count_24__N_543_adj_1404[19]), 
           .\count_24__N_543[20] (count_24__N_543_adj_1404[20]), .\count2[17] (count2[17]), 
           .\count2[18] (count2[18]), .\count_24__N_543[17] (count_24__N_543_adj_1404[17]), 
           .\count_24__N_543[18] (count_24__N_543_adj_1404[18]), .\count2[15] (count2[15]), 
           .\count2[16] (count2[16]), .\count_24__N_543[15] (count_24__N_543_adj_1404[15]), 
           .\count_24__N_543[16] (count_24__N_543_adj_1404[16]), .\count2[14] (count2[14]), 
           .\count_24__N_543[13] (count_24__N_543_adj_1404[13]), .\count_24__N_543[14] (count_24__N_543_adj_1404[14]), 
           .\count_24__N_543[11] (count_24__N_543_adj_1404[11]), .\count_24__N_543[12] (count_24__N_543_adj_1404[12]), 
           .\count_24__N_543[9] (count_24__N_543_adj_1404[9]), .\count_24__N_543[10] (count_24__N_543_adj_1404[10]), 
           .\count_24__N_543[7] (count_24__N_543_adj_1404[7]), .\count_24__N_543[8] (count_24__N_543_adj_1404[8]), 
           .n18757(n18757), .\fcw_r[6] (fcw_r[6]), .n18785(n18785), .n18705(n18705), 
           .n18717(n18717), .n19839(n19839), .\yinjie_box[1] (yinjie_box[1]), 
           .n18716(n18716), .\count2[1] (count2[1]), .pwm_out2_N_125(pwm_out2_N_125), 
           .n49(n52_adj_1405[1]), .n48(n52_adj_1405[2]), .n47(n52_adj_1405[3]), 
           .n46(n52_adj_1405[4]), .n45(n52_adj_1405[5]), .n44(n52_adj_1405[6]), 
           .n43(n52_adj_1405[7]), .n42(n52_adj_1405[8]), .n41(n52_adj_1405[9]), 
           .n40(n52_adj_1405[10]), .n39(n52_adj_1405[11]), .n38(n52_adj_1405[12]), 
           .n37(n52_adj_1405[13]), .n36(n52_adj_1405[14]), .n35(n52_adj_1405[15]), 
           .n34(n52_adj_1405[16]), .n33(n52_adj_1405[17]), .n32(n52_adj_1405[18]), 
           .n31(n52_adj_1405[19]), .n30(n52_adj_1405[20]), .n29(n52_adj_1405[21]), 
           .n28(n52_adj_1405[22]), .n27(n52_adj_1405[23]), .n26(n52_adj_1405[24]), 
           .\count_24__N_543[5] (count_24__N_543_adj_1404[5]), .\count_24__N_543[6] (count_24__N_543_adj_1404[6]), 
           .\count_24__N_543[3] (count_24__N_543_adj_1404[3]), .\count_24__N_543[4] (count_24__N_543_adj_1404[4]), 
           .\count_24__N_543[2] (count_24__N_543_adj_1404[2]), .n18608(n18608), 
           .n7920(n7919[7])) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(58[5] 67[3])
    DDS_U7 u_DDS_1 (.n19846(n19846), .\fcw_r[0] (fcw_r_adj_1408[0]), .clk_N_168(clk_N_168), 
           .n18785(n18785), .\count1[24] (count1[24]), .GND_net(GND_net), 
           .n106(n105[24]), .\count1[22] (count1[22]), .\count1[23] (count1[23]), 
           .n108(n105[22]), .n107(n105[23]), .\count1[20] (count1[20]), 
           .\count1[21] (count1[21]), .n110(n105[20]), .n109(n105[21]), 
           .\count1[18] (count1[18]), .\count1[19] (count1[19]), .n112(n105[18]), 
           .n111(n105[19]), .\count1[16] (count1[16]), .\count1[17] (count1[17]), 
           .n114(n105[16]), .n113(n105[17]), .\count1[14] (count1[14]), 
           .\count1[15] (count1[15]), .n116(n105[14]), .n115(n105[15]), 
           .n118(n105[12]), .n117(n105[13]), .\fcw_r[10] (fcw_r_adj_1408[10]), 
           .n120(n105[10]), .n119(n105[11]), .\fcw_r[8] (fcw_r_adj_1408[8]), 
           .\fcw_r[9] (fcw_r_adj_1408[9]), .n122(n105[8]), .n121(n105[9]), 
           .\fcw_r[6] (fcw_r_adj_1408[6]), .\fcw_r[7] (fcw_r_adj_1408[7]), 
           .n124(n105[6]), .n123(n105[7]), .\fcw_r[4] (fcw_r_adj_1408[4]), 
           .\fcw_r[5] (fcw_r_adj_1408[5]), .n126(n105[4]), .n125(n105[5]), 
           .\fcw_r[2] (fcw_r_adj_1408[2]), .\fcw_r[3] (fcw_r_adj_1408[3]), 
           .n128(n105[2]), .n127(n105[3]), .n25(n184[0]), .\fcw_r[1] (fcw_r_adj_1408[1]), 
           .n129(n105[1]), .yinjie({yinjie}), .\yinjie_box[1] (yinjie_box[1]), 
           .\fcw_r_15__N_527[0] (fcw_r_15__N_527[0]), .pwm_out2_N_125(pwm_out2_N_125), 
           .n132({n132}), .stat(stat), .\fcw_r_15__N_495[8] (fcw_r_15__N_495[8]), 
           .clk__inv(clk__inv)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(47[5] 56[3])
    DDS_U8 u_DDS_13 (.\count13[23] (count13[23]), .GND_net(GND_net), .\count13[24] (count13[24]), 
           .\count_24__N_543[23] (count_24__N_543_adj_1406[23]), .\count_24__N_543[24] (count_24__N_543_adj_1406[24]), 
           .\count13[21] (count13[21]), .\count13[22] (count13[22]), .\count_24__N_543[21] (count_24__N_543_adj_1406[21]), 
           .\count_24__N_543[22] (count_24__N_543_adj_1406[22]), .\count13[19] (count13[19]), 
           .\count13[20] (count13[20]), .\count_24__N_543[19] (count_24__N_543_adj_1406[19]), 
           .\count_24__N_543[20] (count_24__N_543_adj_1406[20]), .\count13[17] (count13[17]), 
           .\count13[18] (count13[18]), .\count_24__N_543[17] (count_24__N_543_adj_1406[17]), 
           .\count_24__N_543[18] (count_24__N_543_adj_1406[18]), .\count13[15] (count13[15]), 
           .\count13[16] (count13[16]), .\count_24__N_543[15] (count_24__N_543_adj_1406[15]), 
           .\count_24__N_543[16] (count_24__N_543_adj_1406[16]), .\count13[14] (count13[14]), 
           .\count_24__N_543[13] (count_24__N_543_adj_1406[13]), .\count_24__N_543[14] (count_24__N_543_adj_1406[14]), 
           .\fcw_r[10] (fcw_r_adj_1408[10]), .\count_24__N_543[11] (count_24__N_543_adj_1406[11]), 
           .\count_24__N_543[12] (count_24__N_543_adj_1406[12]), .\fcw_r[8] (fcw_r_adj_1408[8]), 
           .\fcw_r[9] (fcw_r_adj_1408[9]), .\count_24__N_543[9] (count_24__N_543_adj_1406[9]), 
           .\count_24__N_543[10] (count_24__N_543_adj_1406[10]), .\fcw_r[6] (fcw_r_adj_1408[6]), 
           .\fcw_r[7] (fcw_r_adj_1408[7]), .\count_24__N_543[7] (count_24__N_543_adj_1406[7]), 
           .\count_24__N_543[8] (count_24__N_543_adj_1406[8]), .\fcw_r[4] (fcw_r_adj_1408[4]), 
           .\fcw_r[5] (fcw_r_adj_1408[5]), .\count_24__N_543[5] (count_24__N_543_adj_1406[5]), 
           .\count_24__N_543[6] (count_24__N_543_adj_1406[6]), .\fcw_r[2] (fcw_r_adj_1408[2]), 
           .\fcw_r[3] (fcw_r_adj_1408[3]), .\count_24__N_543[3] (count_24__N_543_adj_1406[3]), 
           .\count_24__N_543[4] (count_24__N_543_adj_1406[4]), .\count13[1] (count13[1]), 
           .\fcw_r[0] (fcw_r_adj_1408[0]), .\fcw_r[1] (fcw_r_adj_1408[1]), 
           .\count_24__N_543[2] (count_24__N_543_adj_1406[2]), .clk(clk), 
           .clk__inv(clk__inv), .rst_n_c(rst_n_c), .key_pa_c(key_pa_c), 
           .pwm_out2_N_125(pwm_out2_N_125), .clk_N_168(clk_N_168), .n49(n52_adj_1407[1]), 
           .n48(n52_adj_1407[2]), .n47(n52_adj_1407[3]), .n46(n52_adj_1407[4]), 
           .n45(n52_adj_1407[5]), .n44(n52_adj_1407[6]), .n43(n52_adj_1407[7]), 
           .n42(n52_adj_1407[8]), .n41(n52_adj_1407[9]), .n40(n52_adj_1407[10]), 
           .n39(n52_adj_1407[11]), .n38(n52_adj_1407[12]), .n37(n52_adj_1407[13]), 
           .n36(n52_adj_1407[14]), .n35(n52_adj_1407[15]), .n34(n52_adj_1407[16]), 
           .n33(n52_adj_1407[17]), .n32(n52_adj_1407[18]), .n31(n52_adj_1407[19]), 
           .n30(n52_adj_1407[20]), .n29(n52_adj_1407[21]), .n28(n52_adj_1407[22]), 
           .n27(n52_adj_1407[23]), .n26(n52_adj_1407[24])) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(179[5] 188[3])
    DDS_U9 u_DDS_12 (.\count12[24] (count12[24]), .GND_net(GND_net), .n106(n105_adj_1420[24]), 
           .\count12[22] (count12[22]), .\count12[23] (count12[23]), .n108(n105_adj_1420[22]), 
           .n107(n105_adj_1420[23]), .\count12[20] (count12[20]), .\count12[21] (count12[21]), 
           .n110(n105_adj_1420[20]), .n109(n105_adj_1420[21]), .\count12[18] (count12[18]), 
           .\count12[19] (count12[19]), .n112(n105_adj_1420[18]), .n111(n105_adj_1420[19]), 
           .\count12[16] (count12[16]), .\count12[17] (count12[17]), .n114(n105_adj_1420[16]), 
           .n113(n105_adj_1420[17]), .\count12[14] (count12[14]), .\count12[15] (count12[15]), 
           .n116(n105_adj_1420[14]), .n115(n105_adj_1420[15]), .n118(n105_adj_1420[12]), 
           .n117(n105_adj_1420[13]), .\fcw_r[2] (fcw_r_adj_1433[2]), .n120(n105_adj_1420[10]), 
           .n119(n105_adj_1420[11]), .\fcw_r[0] (fcw_r_adj_1412[0]), .\fcw_r[1] (fcw_r_adj_1433[1]), 
           .n122(n105_adj_1420[8]), .n121(n105_adj_1420[9]), .n124(n105_adj_1420[6]), 
           .n123(n105_adj_1420[7]), .n126(n105_adj_1420[4]), .n125(n105_adj_1420[5]), 
           .n128(n105_adj_1420[2]), .n127(n105_adj_1420[3]), .n25(n184_adj_1422[0]), 
           .n129(n105_adj_1420[1]), .clk_N_168(clk_N_168), .pwm_out2_N_125(pwm_out2_N_125), 
           .n132({n132_adj_1421}), .n18757(n18757), .\fcw_r_15__N_495[11] (\fcw_r_15__N_495[11] ), 
           .yinjie({yinjie}), .n18785(n18785), .n18784(n18784), .n19846(n19846), 
           .\yinjie_box[1] (yinjie_box[1]), .\fcw_r_15__N_527[0] (fcw_r_15__N_527[0])) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(168[5] 177[3])
    DDS_U10 u_DDS_11 (.clk_N_168(clk_N_168), .n18705(n18705), .\count11[23] (count11[23]), 
            .GND_net(GND_net), .\count11[24] (count11[24]), .\count_24__N_543[23] (count_24__N_543_adj_1400[23]), 
            .\count_24__N_543[24] (count_24__N_543_adj_1400[24]), .\count11[21] (count11[21]), 
            .\count11[22] (count11[22]), .\count_24__N_543[21] (count_24__N_543_adj_1400[21]), 
            .\count_24__N_543[22] (count_24__N_543_adj_1400[22]), .\count11[19] (count11[19]), 
            .\count11[20] (count11[20]), .\count_24__N_543[19] (count_24__N_543_adj_1400[19]), 
            .\count_24__N_543[20] (count_24__N_543_adj_1400[20]), .\count11[17] (count11[17]), 
            .\count11[18] (count11[18]), .\count_24__N_543[17] (count_24__N_543_adj_1400[17]), 
            .\count_24__N_543[18] (count_24__N_543_adj_1400[18]), .\count11[15] (count11[15]), 
            .\count11[16] (count11[16]), .\count_24__N_543[15] (count_24__N_543_adj_1400[15]), 
            .\count_24__N_543[16] (count_24__N_543_adj_1400[16]), .\count11[14] (count11[14]), 
            .\count_24__N_543[13] (count_24__N_543_adj_1400[13]), .\count_24__N_543[14] (count_24__N_543_adj_1400[14]), 
            .\count_24__N_543[11] (count_24__N_543_adj_1400[11]), .\count_24__N_543[12] (count_24__N_543_adj_1400[12]), 
            .\count_24__N_543[9] (count_24__N_543_adj_1400[9]), .\count_24__N_543[10] (count_24__N_543_adj_1400[10]), 
            .\count_24__N_543[7] (count_24__N_543_adj_1400[7]), .\count_24__N_543[8] (count_24__N_543_adj_1400[8]), 
            .\fcw_r[6] (fcw_r_adj_1425[6]), .\count_24__N_543[5] (count_24__N_543_adj_1400[5]), 
            .\count_24__N_543[6] (count_24__N_543_adj_1400[6]), .\count_24__N_543[3] (count_24__N_543_adj_1400[3]), 
            .\count_24__N_543[4] (count_24__N_543_adj_1400[4]), .\count11[1] (count11[1]), 
            .\count_24__N_543[2] (count_24__N_543_adj_1400[2]), .n18757(n18757), 
            .n18716(n18716), .\fcw_r_15__N_495[11] (\fcw_r_15__N_495[11] ), 
            .n18634(n18634), .n18608(n18608), .pwm_out2_N_125(pwm_out2_N_125), 
            .n49(n52_adj_1401[1]), .n48(n52_adj_1401[2]), .n47(n52_adj_1401[3]), 
            .n46(n52_adj_1401[4]), .n45(n52_adj_1401[5]), .n44(n52_adj_1401[6]), 
            .n43(n52_adj_1401[7]), .n42(n52_adj_1401[8]), .n41(n52_adj_1401[9]), 
            .n40(n52_adj_1401[10]), .n39(n52_adj_1401[11]), .n38(n52_adj_1401[12]), 
            .n37(n52_adj_1401[13]), .n36(n52_adj_1401[14]), .n35(n52_adj_1401[15]), 
            .n34(n52_adj_1401[16]), .n33(n52_adj_1401[17]), .n32(n52_adj_1401[18]), 
            .n31(n52_adj_1401[19]), .n30(n52_adj_1401[20]), .n29(n52_adj_1401[21]), 
            .n28(n52_adj_1401[22]), .n27(n52_adj_1401[23]), .n26(n52_adj_1401[24]), 
            .n18717(n18717), .n19839(n19839), .n19840(n19840), .n18785(n18785), 
            .n18784(n18784), .\fcw_r_15__N_495[8] (fcw_r_15__N_495[8]), 
            .\fcw_r_15__N_495[9] (\fcw_r_15__N_495[9] ), .\fcw_r_15__N_495[10] (\fcw_r_15__N_495[10] )) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(157[5] 166[3])
    DDS_U11 u_DDS_10 (.\fcw_r[2] (fcw_r_adj_1426[2]), .clk_N_168(clk_N_168), 
            .n18785(n18785), .\count10[24] (count10[24]), .GND_net(GND_net), 
            .\count_24__N_543[24] (count_24__N_543_adj_1423[24]), .\count10[22] (count10[22]), 
            .\count10[23] (count10[23]), .\count_24__N_543[22] (count_24__N_543_adj_1423[22]), 
            .\count_24__N_543[23] (count_24__N_543_adj_1423[23]), .\count10[20] (count10[20]), 
            .\count10[21] (count10[21]), .\count_24__N_543[20] (count_24__N_543_adj_1423[20]), 
            .\count_24__N_543[21] (count_24__N_543_adj_1423[21]), .\count10[18] (count10[18]), 
            .\count10[19] (count10[19]), .\count_24__N_543[18] (count_24__N_543_adj_1423[18]), 
            .\count_24__N_543[19] (count_24__N_543_adj_1423[19]), .\count10[16] (count10[16]), 
            .\count10[17] (count10[17]), .\count_24__N_543[16] (count_24__N_543_adj_1423[16]), 
            .\count_24__N_543[17] (count_24__N_543_adj_1423[17]), .\count10[14] (count10[14]), 
            .\count10[15] (count10[15]), .\count_24__N_543[14] (count_24__N_543_adj_1423[14]), 
            .\count_24__N_543[15] (count_24__N_543_adj_1423[15]), .\count_24__N_543[12] (count_24__N_543_adj_1423[12]), 
            .\count_24__N_543[13] (count_24__N_543_adj_1423[13]), .\count_24__N_543[10] (count_24__N_543_adj_1423[10]), 
            .\count_24__N_543[11] (count_24__N_543_adj_1423[11]), .\count_24__N_543[8] (count_24__N_543_adj_1423[8]), 
            .\count_24__N_543[9] (count_24__N_543_adj_1423[9]), .\count_24__N_543[6] (count_24__N_543_adj_1423[6]), 
            .\count_24__N_543[7] (count_24__N_543_adj_1423[7]), .\count_24__N_543[4] (count_24__N_543_adj_1423[4]), 
            .\count_24__N_543[5] (count_24__N_543_adj_1423[5]), .\count10[2] (count10[2]), 
            .\count_24__N_543[3] (count_24__N_543_adj_1423[3]), .pwm_out2_N_125(pwm_out2_N_125), 
            .n48(n52_adj_1424[2]), .n47(n52_adj_1424[3]), .n46(n52_adj_1424[4]), 
            .n45(n52_adj_1424[5]), .n44(n52_adj_1424[6]), .n43(n52_adj_1424[7]), 
            .n42(n52_adj_1424[8]), .n41(n52_adj_1424[9]), .n40(n52_adj_1424[10]), 
            .n39(n52_adj_1424[11]), .n38(n52_adj_1424[12]), .n37(n52_adj_1424[13]), 
            .n36(n52_adj_1424[14]), .n35(n52_adj_1424[15]), .n34(n52_adj_1424[16]), 
            .n33(n52_adj_1424[17]), .n32(n52_adj_1424[18]), .n31(n52_adj_1424[19]), 
            .n30(n52_adj_1424[20]), .n29(n52_adj_1424[21]), .n28(n52_adj_1424[22]), 
            .n27(n52_adj_1424[23]), .n26(n52_adj_1424[24]), .n18784(n18784), 
            .\fcw_r_15__N_495[8] (fcw_r_15__N_495[8]), .\fcw_r_15__N_495[5] (\fcw_r_15__N_495[5] ), 
            .\fcw_r_15__N_495[6] (\fcw_r_15__N_495[6] ), .\fcw_r_15__N_495[8]_adj_10 (\fcw_r_15__N_495[8] ), 
            .\fcw_r_15__N_495[9] (\fcw_r_15__N_495[9] ), .\fcw_r_15__N_495[10] (\fcw_r_15__N_495[10] ), 
            .n19846(n19846), .\yinjie[2] (yinjie[2]), .n18757(n18757), 
            .\fcw_r_15__N_495[11] (\fcw_r_15__N_495[11] ), .n18716(n18716), 
            .n18634(n18634), .n15966(n15966), .n18690(n18690), .n18705(n18705), 
            .n16936(n16936), .n10972(n10972)) /* synthesis syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(146[5] 155[3])
    sin_rom sin2 (.\u_count2[24] (u_count2[24]), .\u_count2[23] (u_count2[23]), 
            .\u_count2[22] (u_count2[22]), .\u_count2[21] (u_count2[21]), 
            .\u_count2[20] (u_count2[20]), .\u_count2[19] (u_count2[19]), 
            .\u_count2[18] (u_count2[18]), .\u_count2[17] (u_count2[17]), 
            .\u_count2[16] (u_count2[16]), .\u_count2[15] (u_count2[15]), 
            .\u_count2[14] (u_count2[14]), .clk(clk), .\en[1] (en[1]), 
            .GND_net(GND_net), .data_out2({data_out2[11:1], \data_out2[0] }), 
            .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(38[10] 44[4])
    sin_rom_U12 sin1 (.\u_count1[24] (u_count1[24]), .\u_count1[23] (u_count1[23]), 
            .\u_count1[22] (u_count1[22]), .\u_count1[21] (u_count1[21]), 
            .\u_count1[20] (u_count1[20]), .\u_count1[19] (u_count1[19]), 
            .\u_count1[18] (u_count1[18]), .\u_count1[17] (u_count1[17]), 
            .\u_count1[16] (u_count1[16]), .\u_count1[15] (u_count1[15]), 
            .\u_count1[14] (u_count1[14]), .clk(clk), .\en[0] (en[0]), 
            .GND_net(GND_net), .data_out1({data_out1[11:1], \data_out1[0] }), 
            .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(31[10] 37[4])
    
endmodule
//
// Verilog Description of module DDS
//

module DDS (\fcw_r[8] , clk_N_168, n18785, \count9[23] , GND_net, 
            \count9[24] , \count_24__N_543[23] , \count_24__N_543[24] , 
            \count9[21] , \count9[22] , \count_24__N_543[21] , \count_24__N_543[22] , 
            \count9[19] , \count9[20] , \count_24__N_543[19] , \count_24__N_543[20] , 
            \count9[17] , \count9[18] , \count_24__N_543[17] , \count_24__N_543[18] , 
            \count9[15] , \count9[16] , \count_24__N_543[15] , \count_24__N_543[16] , 
            \count9[14] , \count_24__N_543[13] , \count_24__N_543[14] , 
            \count_24__N_543[11] , \count_24__N_543[12] , \count_24__N_543[9] , 
            \count_24__N_543[10] , \count_24__N_543[7] , \count_24__N_543[8] , 
            \count_24__N_543[5] , \count_24__N_543[6] , \count_24__N_543[3] , 
            \count_24__N_543[4] , \count9[1] , \count_24__N_543[2] , pwm_out2_N_125, 
            n49, n48, n47, n46, n45, n44, n43, n42, n41, n40, 
            n39, n38, n37, n36, n35, n34, n33, n32, n31, n30, 
            n29, n28, n27, n26, n18784, n18757) /* synthesis syn_module_defined=1 */ ;
    output \fcw_r[8] ;
    input clk_N_168;
    input n18785;
    output \count9[23] ;
    input GND_net;
    output \count9[24] ;
    output \count_24__N_543[23] ;
    output \count_24__N_543[24] ;
    output \count9[21] ;
    output \count9[22] ;
    output \count_24__N_543[21] ;
    output \count_24__N_543[22] ;
    output \count9[19] ;
    output \count9[20] ;
    output \count_24__N_543[19] ;
    output \count_24__N_543[20] ;
    output \count9[17] ;
    output \count9[18] ;
    output \count_24__N_543[17] ;
    output \count_24__N_543[18] ;
    output \count9[15] ;
    output \count9[16] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[16] ;
    output \count9[14] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[14] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[12] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[10] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[8] ;
    output \count_24__N_543[5] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[3] ;
    output \count_24__N_543[4] ;
    output \count9[1] ;
    output \count_24__N_543[2] ;
    input pwm_out2_N_125;
    input n49;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    input n18784;
    input n18757;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15429, n15428, n15427, n15426, n15425, n15424;
    wire [24:0]count9;   // d:/fpga_project/lattice_diamond/piano/speaker.v(13[52:58])
    
    wire n15423, n15422;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15421, n15420, n15419;
    
    FD1S3AX fcw_r_i1 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[8] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D add_2212_24 (.A0(\count9[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count9[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15429), .S0(\count_24__N_543[23] ), .S1(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_24.INIT0 = 16'h5aaa;
    defparam add_2212_24.INIT1 = 16'h5aaa;
    defparam add_2212_24.INJECT1_0 = "NO";
    defparam add_2212_24.INJECT1_1 = "NO";
    CCU2D add_2212_22 (.A0(\count9[21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count9[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15428), .COUT(n15429), .S0(\count_24__N_543[21] ), 
          .S1(\count_24__N_543[22] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_22.INIT0 = 16'h5aaa;
    defparam add_2212_22.INIT1 = 16'h5aaa;
    defparam add_2212_22.INJECT1_0 = "NO";
    defparam add_2212_22.INJECT1_1 = "NO";
    CCU2D add_2212_20 (.A0(\count9[19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count9[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15427), .COUT(n15428), .S0(\count_24__N_543[19] ), 
          .S1(\count_24__N_543[20] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_20.INIT0 = 16'h5aaa;
    defparam add_2212_20.INIT1 = 16'h5aaa;
    defparam add_2212_20.INJECT1_0 = "NO";
    defparam add_2212_20.INJECT1_1 = "NO";
    CCU2D add_2212_18 (.A0(\count9[17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count9[18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15426), .COUT(n15427), .S0(\count_24__N_543[17] ), 
          .S1(\count_24__N_543[18] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_18.INIT0 = 16'h5aaa;
    defparam add_2212_18.INIT1 = 16'h5aaa;
    defparam add_2212_18.INJECT1_0 = "NO";
    defparam add_2212_18.INJECT1_1 = "NO";
    CCU2D add_2212_16 (.A0(\count9[15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count9[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15425), .COUT(n15426), .S0(\count_24__N_543[15] ), 
          .S1(\count_24__N_543[16] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_16.INIT0 = 16'h5aaa;
    defparam add_2212_16.INIT1 = 16'h5aaa;
    defparam add_2212_16.INJECT1_0 = "NO";
    defparam add_2212_16.INJECT1_1 = "NO";
    CCU2D add_2212_14 (.A0(count9[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count9[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15424), .COUT(n15425), .S0(\count_24__N_543[13] ), .S1(\count_24__N_543[14] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_14.INIT0 = 16'h5aaa;
    defparam add_2212_14.INIT1 = 16'h5aaa;
    defparam add_2212_14.INJECT1_0 = "NO";
    defparam add_2212_14.INJECT1_1 = "NO";
    CCU2D add_2212_12 (.A0(count9[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count9[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15423), .COUT(n15424), .S0(\count_24__N_543[11] ), .S1(\count_24__N_543[12] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_12.INIT0 = 16'h5aaa;
    defparam add_2212_12.INIT1 = 16'h5aaa;
    defparam add_2212_12.INJECT1_0 = "NO";
    defparam add_2212_12.INJECT1_1 = "NO";
    CCU2D add_2212_10 (.A0(count9[9]), .B0(fcw_r[9]), .C0(GND_net), .D0(GND_net), 
          .A1(count9[10]), .B1(fcw_r[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15422), .COUT(n15423), .S0(\count_24__N_543[9] ), .S1(\count_24__N_543[10] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_10.INIT0 = 16'h5666;
    defparam add_2212_10.INIT1 = 16'h5666;
    defparam add_2212_10.INJECT1_0 = "NO";
    defparam add_2212_10.INJECT1_1 = "NO";
    CCU2D add_2212_8 (.A0(count9[7]), .B0(fcw_r[10]), .C0(GND_net), .D0(GND_net), 
          .A1(count9[8]), .B1(\fcw_r[8] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15421), .COUT(n15422), .S0(\count_24__N_543[7] ), .S1(\count_24__N_543[8] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_8.INIT0 = 16'h5666;
    defparam add_2212_8.INIT1 = 16'h5666;
    defparam add_2212_8.INJECT1_0 = "NO";
    defparam add_2212_8.INJECT1_1 = "NO";
    CCU2D add_2212_6 (.A0(count9[5]), .B0(\fcw_r[8] ), .C0(GND_net), .D0(GND_net), 
          .A1(count9[6]), .B1(fcw_r[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15420), .COUT(n15421), .S0(\count_24__N_543[5] ), .S1(\count_24__N_543[6] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_6.INIT0 = 16'h5666;
    defparam add_2212_6.INIT1 = 16'h5666;
    defparam add_2212_6.INJECT1_0 = "NO";
    defparam add_2212_6.INJECT1_1 = "NO";
    CCU2D add_2212_4 (.A0(count9[3]), .B0(fcw_r[10]), .C0(GND_net), .D0(GND_net), 
          .A1(count9[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15419), .COUT(n15420), .S0(\count_24__N_543[3] ), .S1(\count_24__N_543[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_4.INIT0 = 16'h5666;
    defparam add_2212_4.INIT1 = 16'h5aaa;
    defparam add_2212_4.INJECT1_0 = "NO";
    defparam add_2212_4.INJECT1_1 = "NO";
    CCU2D add_2212_2 (.A0(\count9[1] ), .B0(\fcw_r[8] ), .C0(GND_net), 
          .D0(GND_net), .A1(count9[2]), .B1(fcw_r[9]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15419), .S1(\count_24__N_543[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2212_2.INIT0 = 16'h7000;
    defparam add_2212_2.INIT1 = 16'h5666;
    defparam add_2212_2.INJECT1_0 = "NO";
    defparam add_2212_2.INJECT1_1 = "NO";
    FD1S3DX count__i1 (.D(n49), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count9[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i1.GSR = "DISABLED";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count9[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count9[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count9[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count9[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count9[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count9[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    FD1S3AX fcw_r_i2 (.D(n18784), .CK(clk_N_168), .Q(fcw_r[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(n18757), .CK(clk_N_168), .Q(fcw_r[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=135, LSE_RLINE=144 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U0
//

module DDS_U0 (\fcw_r[8] , clk_N_168, n18785, \count8[23] , GND_net, 
            \count8[24] , \count_24__N_543[23] , \count_24__N_543[24] , 
            \count8[21] , \count8[22] , \count_24__N_543[21] , \count_24__N_543[22] , 
            \count8[19] , \count8[20] , \count_24__N_543[19] , \count_24__N_543[20] , 
            \count8[17] , \count8[18] , \count_24__N_543[17] , \count_24__N_543[18] , 
            \count8[15] , \count8[16] , \count_24__N_543[15] , \count_24__N_543[16] , 
            \count8[14] , \count_24__N_543[13] , \count_24__N_543[14] , 
            \count_24__N_543[11] , \count_24__N_543[12] , \count_24__N_543[9] , 
            \count_24__N_543[10] , \count_24__N_543[7] , \count_24__N_543[8] , 
            \count_24__N_543[5] , \count_24__N_543[6] , \count_24__N_543[3] , 
            \count_24__N_543[4] , \count8[1] , \count_24__N_543[2] , pwm_out2_N_125, 
            n49, n48, n47, n46, n45, n44, n43, n42, n41, n40, 
            n39, n38, n37, n36, n35, n34, n33, n32, n31, n30, 
            n29, n28, n27, n26, n18784, n18757) /* synthesis syn_module_defined=1 */ ;
    output \fcw_r[8] ;
    input clk_N_168;
    input n18785;
    output \count8[23] ;
    input GND_net;
    output \count8[24] ;
    output \count_24__N_543[23] ;
    output \count_24__N_543[24] ;
    output \count8[21] ;
    output \count8[22] ;
    output \count_24__N_543[21] ;
    output \count_24__N_543[22] ;
    output \count8[19] ;
    output \count8[20] ;
    output \count_24__N_543[19] ;
    output \count_24__N_543[20] ;
    output \count8[17] ;
    output \count8[18] ;
    output \count_24__N_543[17] ;
    output \count_24__N_543[18] ;
    output \count8[15] ;
    output \count8[16] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[16] ;
    output \count8[14] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[14] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[12] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[10] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[8] ;
    output \count_24__N_543[5] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[3] ;
    output \count_24__N_543[4] ;
    output \count8[1] ;
    output \count_24__N_543[2] ;
    input pwm_out2_N_125;
    input n49;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    input n18784;
    input n18757;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15416, n15415, n15414, n15413, n15412, n15411;
    wire [24:0]count8;   // d:/fpga_project/lattice_diamond/piano/speaker.v(13[33:39])
    
    wire n15410, n15409;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15408, n15407, n15406;
    
    FD1S3AX fcw_r_i1 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[8] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D add_2211_24 (.A0(\count8[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count8[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15416), .S0(\count_24__N_543[23] ), .S1(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_24.INIT0 = 16'h5aaa;
    defparam add_2211_24.INIT1 = 16'h5aaa;
    defparam add_2211_24.INJECT1_0 = "NO";
    defparam add_2211_24.INJECT1_1 = "NO";
    CCU2D add_2211_22 (.A0(\count8[21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count8[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15415), .COUT(n15416), .S0(\count_24__N_543[21] ), 
          .S1(\count_24__N_543[22] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_22.INIT0 = 16'h5aaa;
    defparam add_2211_22.INIT1 = 16'h5aaa;
    defparam add_2211_22.INJECT1_0 = "NO";
    defparam add_2211_22.INJECT1_1 = "NO";
    CCU2D add_2211_20 (.A0(\count8[19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count8[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15414), .COUT(n15415), .S0(\count_24__N_543[19] ), 
          .S1(\count_24__N_543[20] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_20.INIT0 = 16'h5aaa;
    defparam add_2211_20.INIT1 = 16'h5aaa;
    defparam add_2211_20.INJECT1_0 = "NO";
    defparam add_2211_20.INJECT1_1 = "NO";
    CCU2D add_2211_18 (.A0(\count8[17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count8[18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15413), .COUT(n15414), .S0(\count_24__N_543[17] ), 
          .S1(\count_24__N_543[18] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_18.INIT0 = 16'h5aaa;
    defparam add_2211_18.INIT1 = 16'h5aaa;
    defparam add_2211_18.INJECT1_0 = "NO";
    defparam add_2211_18.INJECT1_1 = "NO";
    CCU2D add_2211_16 (.A0(\count8[15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count8[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15412), .COUT(n15413), .S0(\count_24__N_543[15] ), 
          .S1(\count_24__N_543[16] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_16.INIT0 = 16'h5aaa;
    defparam add_2211_16.INIT1 = 16'h5aaa;
    defparam add_2211_16.INJECT1_0 = "NO";
    defparam add_2211_16.INJECT1_1 = "NO";
    CCU2D add_2211_14 (.A0(count8[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count8[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15411), .COUT(n15412), .S0(\count_24__N_543[13] ), .S1(\count_24__N_543[14] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_14.INIT0 = 16'h5aaa;
    defparam add_2211_14.INIT1 = 16'h5aaa;
    defparam add_2211_14.INJECT1_0 = "NO";
    defparam add_2211_14.INJECT1_1 = "NO";
    CCU2D add_2211_12 (.A0(count8[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count8[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15410), .COUT(n15411), .S0(\count_24__N_543[11] ), .S1(\count_24__N_543[12] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_12.INIT0 = 16'h5aaa;
    defparam add_2211_12.INIT1 = 16'h5aaa;
    defparam add_2211_12.INJECT1_0 = "NO";
    defparam add_2211_12.INJECT1_1 = "NO";
    CCU2D add_2211_10 (.A0(count8[9]), .B0(fcw_r[9]), .C0(GND_net), .D0(GND_net), 
          .A1(count8[10]), .B1(fcw_r[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15409), .COUT(n15410), .S0(\count_24__N_543[9] ), .S1(\count_24__N_543[10] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_10.INIT0 = 16'h5666;
    defparam add_2211_10.INIT1 = 16'h5666;
    defparam add_2211_10.INJECT1_0 = "NO";
    defparam add_2211_10.INJECT1_1 = "NO";
    CCU2D add_2211_8 (.A0(count8[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count8[8]), .B1(\fcw_r[8] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15408), .COUT(n15409), .S0(\count_24__N_543[7] ), .S1(\count_24__N_543[8] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_8.INIT0 = 16'h5aaa;
    defparam add_2211_8.INIT1 = 16'h5666;
    defparam add_2211_8.INJECT1_0 = "NO";
    defparam add_2211_8.INJECT1_1 = "NO";
    CCU2D add_2211_6 (.A0(count8[5]), .B0(fcw_r[9]), .C0(GND_net), .D0(GND_net), 
          .A1(count8[6]), .B1(fcw_r[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15407), .COUT(n15408), .S0(\count_24__N_543[5] ), .S1(\count_24__N_543[6] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_6.INIT0 = 16'h5666;
    defparam add_2211_6.INIT1 = 16'h5666;
    defparam add_2211_6.INJECT1_0 = "NO";
    defparam add_2211_6.INJECT1_1 = "NO";
    CCU2D add_2211_4 (.A0(count8[3]), .B0(fcw_r[10]), .C0(GND_net), .D0(GND_net), 
          .A1(count8[4]), .B1(\fcw_r[8] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15406), .COUT(n15407), .S0(\count_24__N_543[3] ), .S1(\count_24__N_543[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_4.INIT0 = 16'h5666;
    defparam add_2211_4.INIT1 = 16'h5666;
    defparam add_2211_4.INJECT1_0 = "NO";
    defparam add_2211_4.INJECT1_1 = "NO";
    CCU2D add_2211_2 (.A0(\count8[1] ), .B0(\fcw_r[8] ), .C0(GND_net), 
          .D0(GND_net), .A1(count8[2]), .B1(fcw_r[9]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15406), .S1(\count_24__N_543[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2211_2.INIT0 = 16'h7000;
    defparam add_2211_2.INIT1 = 16'h5666;
    defparam add_2211_2.INJECT1_0 = "NO";
    defparam add_2211_2.INJECT1_1 = "NO";
    FD1S3DX count__i1 (.D(n49), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count8[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i1.GSR = "DISABLED";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count8[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count8[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count8[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count8[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count8[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count8[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    FD1S3AX fcw_r_i2 (.D(n18784), .CK(clk_N_168), .Q(fcw_r[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(n18757), .CK(clk_N_168), .Q(fcw_r[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=124, LSE_RLINE=133 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U1
//

module DDS_U1 (clk_N_168, n18705, \count7[24] , GND_net, n106, \count7[22] , 
            \count7[23] , n108, n107, \count7[20] , \count7[21] , 
            n110, n109, \count7[18] , \count7[19] , n112, n111, 
            \count7[16] , \count7[17] , n114, n113, \count7[14] , 
            \count7[15] , n116, n115, n118, n117, n120, n119, 
            \fcw_r[8] , n122, n121, n124, n123, n126, n125, n128, 
            n127, n25, n129, pwm_out2_N_125, n132, n18717, n19839, 
            n19840, n18785, n18784, n18757) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    input n18705;
    output \count7[24] ;
    input GND_net;
    output n106;
    output \count7[22] ;
    output \count7[23] ;
    output n108;
    output n107;
    output \count7[20] ;
    output \count7[21] ;
    output n110;
    output n109;
    output \count7[18] ;
    output \count7[19] ;
    output n112;
    output n111;
    output \count7[16] ;
    output \count7[17] ;
    output n114;
    output n113;
    output \count7[14] ;
    output \count7[15] ;
    output n116;
    output n115;
    output n118;
    output n117;
    output n120;
    output n119;
    output \fcw_r[8] ;
    output n122;
    output n121;
    output n124;
    output n123;
    output n126;
    output n125;
    output n128;
    output n127;
    output n25;
    output n129;
    input pwm_out2_N_125;
    input [24:0]n132;
    input n18717;
    input n19839;
    input n19840;
    input n18785;
    input n18784;
    input n18757;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15734, n15733, n15732, n15731, n15730, n15729, n15728;
    wire [24:0]n184;
    
    wire n15727, n15726, n15725, n15724, n15723;
    
    FD1S3AX fcw_r_i1 (.D(n18705), .CK(clk_N_168), .Q(fcw_r[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D count_2229_add_4_26 (.A0(\count7[24] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15734), .S0(n106));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_26.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_26.INIT1 = 16'h0000;
    defparam count_2229_add_4_26.INJECT1_0 = "NO";
    defparam count_2229_add_4_26.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_24 (.A0(\count7[22] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count7[23] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15733), .COUT(n15734), .S0(n108), .S1(n107));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_24.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_24.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_24.INJECT1_0 = "NO";
    defparam count_2229_add_4_24.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_22 (.A0(\count7[20] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count7[21] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15732), .COUT(n15733), .S0(n110), .S1(n109));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_22.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_22.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_22.INJECT1_0 = "NO";
    defparam count_2229_add_4_22.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_20 (.A0(\count7[18] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count7[19] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15731), .COUT(n15732), .S0(n112), .S1(n111));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_20.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_20.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_20.INJECT1_0 = "NO";
    defparam count_2229_add_4_20.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_18 (.A0(\count7[16] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count7[17] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15730), .COUT(n15731), .S0(n114), .S1(n113));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_18.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_18.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_18.INJECT1_0 = "NO";
    defparam count_2229_add_4_18.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_16 (.A0(\count7[14] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count7[15] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15729), .COUT(n15730), .S0(n116), .S1(n115));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_16.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_16.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_16.INJECT1_0 = "NO";
    defparam count_2229_add_4_16.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_14 (.A0(n184[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n184[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15728), .COUT(n15729), .S0(n118), .S1(n117));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_14.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_14.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_14.INJECT1_0 = "NO";
    defparam count_2229_add_4_14.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_12 (.A0(fcw_r[10]), .B0(n184[10]), .C0(GND_net), 
          .D0(GND_net), .A1(n184[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15727), .COUT(n15728), .S0(n120), .S1(n119));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_12.INIT0 = 16'h5666;
    defparam count_2229_add_4_12.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_12.INJECT1_0 = "NO";
    defparam count_2229_add_4_12.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_10 (.A0(\fcw_r[8] ), .B0(n184[8]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[9]), .B1(n184[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15726), .COUT(n15727), .S0(n122), .S1(n121));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_10.INIT0 = 16'h5666;
    defparam count_2229_add_4_10.INIT1 = 16'h5666;
    defparam count_2229_add_4_10.INJECT1_0 = "NO";
    defparam count_2229_add_4_10.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_8 (.A0(n184[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n184[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15725), .COUT(n15726), .S0(n124), .S1(n123));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_8.INIT0 = 16'hfaaa;
    defparam count_2229_add_4_8.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_8.INJECT1_0 = "NO";
    defparam count_2229_add_4_8.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_6 (.A0(fcw_r[4]), .B0(n184[4]), .C0(GND_net), 
          .D0(GND_net), .A1(n184[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15724), .COUT(n15725), .S0(n126), .S1(n125));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_6.INIT0 = 16'h5666;
    defparam count_2229_add_4_6.INIT1 = 16'hfaaa;
    defparam count_2229_add_4_6.INJECT1_0 = "NO";
    defparam count_2229_add_4_6.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_4 (.A0(fcw_r[2]), .B0(n184[2]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[3]), .B1(n184[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15723), .COUT(n15724), .S0(n128), .S1(n127));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_4.INIT0 = 16'h5666;
    defparam count_2229_add_4_4.INIT1 = 16'h5666;
    defparam count_2229_add_4_4.INJECT1_0 = "NO";
    defparam count_2229_add_4_4.INJECT1_1 = "NO";
    CCU2D count_2229_add_4_2 (.A0(\fcw_r[8] ), .B0(n25), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[1]), .B1(n184[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n15723), .S1(n129));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229_add_4_2.INIT0 = 16'h7000;
    defparam count_2229_add_4_2.INIT1 = 16'h5666;
    defparam count_2229_add_4_2.INJECT1_0 = "NO";
    defparam count_2229_add_4_2.INJECT1_1 = "NO";
    FD1S3DX count_2229__i0 (.D(n132[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n25)) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i0.GSR = "DISABLED";
    FD1S3AX fcw_r_i2 (.D(n18717), .CK(clk_N_168), .Q(fcw_r[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(n19839), .CK(clk_N_168), .Q(fcw_r[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_i4 (.D(n19840), .CK(clk_N_168), .Q(fcw_r[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_i5 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[8] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_i6 (.D(n18784), .CK(clk_N_168), .Q(fcw_r[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_i7 (.D(n18757), .CK(clk_N_168), .Q(fcw_r[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=113, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i7.GSR = "DISABLED";
    FD1S3DX count_2229__i1 (.D(n132[1]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i1.GSR = "DISABLED";
    FD1S3DX count_2229__i2 (.D(n132[2]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i2.GSR = "DISABLED";
    FD1S3DX count_2229__i3 (.D(n132[3]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i3.GSR = "DISABLED";
    FD1S3DX count_2229__i4 (.D(n132[4]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i4.GSR = "DISABLED";
    FD1S3DX count_2229__i5 (.D(n132[5]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i5.GSR = "DISABLED";
    FD1S3DX count_2229__i6 (.D(n132[6]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i6.GSR = "DISABLED";
    FD1S3DX count_2229__i7 (.D(n132[7]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i7.GSR = "DISABLED";
    FD1S3DX count_2229__i8 (.D(n132[8]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i8.GSR = "DISABLED";
    FD1S3DX count_2229__i9 (.D(n132[9]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i9.GSR = "DISABLED";
    FD1S3DX count_2229__i10 (.D(n132[10]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i10.GSR = "DISABLED";
    FD1S3DX count_2229__i11 (.D(n132[11]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i11.GSR = "DISABLED";
    FD1S3DX count_2229__i12 (.D(n132[12]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i12.GSR = "DISABLED";
    FD1S3DX count_2229__i13 (.D(n132[13]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i13.GSR = "DISABLED";
    FD1S3DX count_2229__i14 (.D(n132[14]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[14] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i14.GSR = "DISABLED";
    FD1S3DX count_2229__i15 (.D(n132[15]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[15] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i15.GSR = "DISABLED";
    FD1S3DX count_2229__i16 (.D(n132[16]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[16] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i16.GSR = "DISABLED";
    FD1S3DX count_2229__i17 (.D(n132[17]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[17] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i17.GSR = "DISABLED";
    FD1S3DX count_2229__i18 (.D(n132[18]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[18] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i18.GSR = "DISABLED";
    FD1S3DX count_2229__i19 (.D(n132[19]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[19] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i19.GSR = "DISABLED";
    FD1S3DX count_2229__i20 (.D(n132[20]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[20] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i20.GSR = "DISABLED";
    FD1S3DX count_2229__i21 (.D(n132[21]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[21] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i21.GSR = "DISABLED";
    FD1S3DX count_2229__i22 (.D(n132[22]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[22] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i22.GSR = "DISABLED";
    FD1S3DX count_2229__i23 (.D(n132[23]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[23] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i23.GSR = "DISABLED";
    FD1S3DX count_2229__i24 (.D(n132[24]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count7[24] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2229__i24.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U2
//

module DDS_U2 (\count6[24] , GND_net, \count_24__N_543[24] , \count6[22] , 
            \count6[23] , \count_24__N_543[22] , \count_24__N_543[23] , 
            \count6[20] , \count6[21] , \count_24__N_543[20] , \count_24__N_543[21] , 
            \count6[18] , \count6[19] , \count_24__N_543[18] , \count_24__N_543[19] , 
            \count6[16] , \count6[17] , \count_24__N_543[16] , \count_24__N_543[17] , 
            \count6[14] , \count6[15] , \count_24__N_543[14] , \count_24__N_543[15] , 
            \count_24__N_543[12] , \count_24__N_543[13] , \fcw_r[2] , 
            \count_24__N_543[10] , \count_24__N_543[11] , \fcw_r[1] , 
            \count_24__N_543[8] , \count_24__N_543[9] , \fcw_r[0] , \count_24__N_543[6] , 
            \count_24__N_543[7] , \fcw_r[4] , \count_24__N_543[4] , \count_24__N_543[5] , 
            \count6[2] , \count_24__N_543[3] , n18717, n18634, \fcw_r_15__N_495[11] , 
            n19839, clk_N_168, pwm_out2_N_125, n48, n47, n46, n45, 
            n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
            n34, n33, n32, n31, n30, n29, n28, n27, n26, \fcw_r_15__N_495[8] , 
            \fcw_r_15__N_495[5] , n16936, n15966, n7920) /* synthesis syn_module_defined=1 */ ;
    output \count6[24] ;
    input GND_net;
    output \count_24__N_543[24] ;
    output \count6[22] ;
    output \count6[23] ;
    output \count_24__N_543[22] ;
    output \count_24__N_543[23] ;
    output \count6[20] ;
    output \count6[21] ;
    output \count_24__N_543[20] ;
    output \count_24__N_543[21] ;
    output \count6[18] ;
    output \count6[19] ;
    output \count_24__N_543[18] ;
    output \count_24__N_543[19] ;
    output \count6[16] ;
    output \count6[17] ;
    output \count_24__N_543[16] ;
    output \count_24__N_543[17] ;
    output \count6[14] ;
    output \count6[15] ;
    output \count_24__N_543[14] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[12] ;
    output \count_24__N_543[13] ;
    input \fcw_r[2] ;
    output \count_24__N_543[10] ;
    output \count_24__N_543[11] ;
    input \fcw_r[1] ;
    output \count_24__N_543[8] ;
    output \count_24__N_543[9] ;
    input \fcw_r[0] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[7] ;
    output \fcw_r[4] ;
    output \count_24__N_543[4] ;
    output \count_24__N_543[5] ;
    output \count6[2] ;
    output \count_24__N_543[3] ;
    input n18717;
    input n18634;
    input \fcw_r_15__N_495[11] ;
    input n19839;
    input clk_N_168;
    input pwm_out2_N_125;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    input \fcw_r_15__N_495[8] ;
    input \fcw_r_15__N_495[5] ;
    input n16936;
    input n15966;
    input n7920;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15404, n15403, n15402, n15401, n15400, n15399, n15398;
    wire [24:0]count6;   // d:/fpga_project/lattice_diamond/piano/speaker.v(12[52:58])
    
    wire n15397, n18694;
    wire [9:0]n6871;
    
    wire n15396, n4, n4_adj_839, n15395;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15394;
    wire [7:0]n7919;
    
    wire n18759;
    
    CCU2D add_15_24 (.A0(\count6[24] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15404), 
          .S0(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_24.INIT0 = 16'h5aaa;
    defparam add_15_24.INIT1 = 16'h0000;
    defparam add_15_24.INJECT1_0 = "NO";
    defparam add_15_24.INJECT1_1 = "NO";
    CCU2D add_15_22 (.A0(\count6[22] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count6[23] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15403), .COUT(n15404), .S0(\count_24__N_543[22] ), .S1(\count_24__N_543[23] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_22.INIT0 = 16'h5aaa;
    defparam add_15_22.INIT1 = 16'h5aaa;
    defparam add_15_22.INJECT1_0 = "NO";
    defparam add_15_22.INJECT1_1 = "NO";
    CCU2D add_15_20 (.A0(\count6[20] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count6[21] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15402), .COUT(n15403), .S0(\count_24__N_543[20] ), .S1(\count_24__N_543[21] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_20.INIT0 = 16'h5aaa;
    defparam add_15_20.INIT1 = 16'h5aaa;
    defparam add_15_20.INJECT1_0 = "NO";
    defparam add_15_20.INJECT1_1 = "NO";
    CCU2D add_15_18 (.A0(\count6[18] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count6[19] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15401), .COUT(n15402), .S0(\count_24__N_543[18] ), .S1(\count_24__N_543[19] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_18.INIT0 = 16'h5aaa;
    defparam add_15_18.INIT1 = 16'h5aaa;
    defparam add_15_18.INJECT1_0 = "NO";
    defparam add_15_18.INJECT1_1 = "NO";
    CCU2D add_15_16 (.A0(\count6[16] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count6[17] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15400), .COUT(n15401), .S0(\count_24__N_543[16] ), .S1(\count_24__N_543[17] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_16.INIT0 = 16'h5aaa;
    defparam add_15_16.INIT1 = 16'h5aaa;
    defparam add_15_16.INJECT1_0 = "NO";
    defparam add_15_16.INJECT1_1 = "NO";
    CCU2D add_15_14 (.A0(\count6[14] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count6[15] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15399), .COUT(n15400), .S0(\count_24__N_543[14] ), .S1(\count_24__N_543[15] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_14.INIT0 = 16'h5aaa;
    defparam add_15_14.INIT1 = 16'h5aaa;
    defparam add_15_14.INJECT1_0 = "NO";
    defparam add_15_14.INJECT1_1 = "NO";
    CCU2D add_15_12 (.A0(count6[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count6[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15398), .COUT(n15399), .S0(\count_24__N_543[12] ), .S1(\count_24__N_543[13] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_12.INIT0 = 16'h5aaa;
    defparam add_15_12.INIT1 = 16'h5aaa;
    defparam add_15_12.INJECT1_0 = "NO";
    defparam add_15_12.INJECT1_1 = "NO";
    CCU2D add_15_10 (.A0(count6[10]), .B0(n18694), .C0(\fcw_r[2] ), .D0(n6871[7]), 
          .A1(count6[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15397), .COUT(n15398), .S0(\count_24__N_543[10] ), .S1(\count_24__N_543[11] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_10.INIT0 = 16'h566a;
    defparam add_15_10.INIT1 = 16'h5aaa;
    defparam add_15_10.INJECT1_0 = "NO";
    defparam add_15_10.INJECT1_1 = "NO";
    CCU2D add_15_8 (.A0(\fcw_r[1] ), .B0(n4), .C0(count6[8]), .D0(GND_net), 
          .A1(\fcw_r[2] ), .B1(n4_adj_839), .C1(count6[9]), .D1(GND_net), 
          .CIN(n15396), .COUT(n15397), .S0(\count_24__N_543[8] ), .S1(\count_24__N_543[9] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_8.INIT0 = 16'h9696;
    defparam add_15_8.INIT1 = 16'h9696;
    defparam add_15_8.INJECT1_0 = "NO";
    defparam add_15_8.INJECT1_1 = "NO";
    CCU2D add_15_6 (.A0(count6[6]), .B0(fcw_r[6]), .C0(GND_net), .D0(GND_net), 
          .A1(n6871[5]), .B1(\fcw_r[0] ), .C1(count6[7]), .D1(GND_net), 
          .CIN(n15395), .COUT(n15396), .S0(\count_24__N_543[6] ), .S1(\count_24__N_543[7] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_6.INIT0 = 16'h5666;
    defparam add_15_6.INIT1 = 16'h9696;
    defparam add_15_6.INJECT1_0 = "NO";
    defparam add_15_6.INJECT1_1 = "NO";
    CCU2D add_15_4 (.A0(count6[4]), .B0(\fcw_r[4] ), .C0(GND_net), .D0(GND_net), 
          .A1(count6[5]), .B1(fcw_r[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15394), .COUT(n15395), .S0(\count_24__N_543[4] ), .S1(\count_24__N_543[5] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_4.INIT0 = 16'h5666;
    defparam add_15_4.INIT1 = 16'h5666;
    defparam add_15_4.INJECT1_0 = "NO";
    defparam add_15_4.INJECT1_1 = "NO";
    CCU2D add_15_2 (.A0(\count6[2] ), .B0(\fcw_r[0] ), .C0(GND_net), .D0(GND_net), 
          .A1(count6[3]), .B1(\fcw_r[1] ), .C1(GND_net), .D1(GND_net), 
          .COUT(n15394), .S1(\count_24__N_543[3] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_2.INIT0 = 16'h7000;
    defparam add_15_2.INIT1 = 16'h5666;
    defparam add_15_2.INJECT1_0 = "NO";
    defparam add_15_2.INJECT1_1 = "NO";
    LUT4 i4148_2_lut_4_lut (.A(n18717), .B(n18634), .C(\fcw_r_15__N_495[11] ), 
         .D(n19839), .Z(n7919[6])) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i4148_2_lut_4_lut.init = 16'h17e8;
    LUT4 i3231_2_lut_rep_577 (.A(n6871[5]), .B(\fcw_r[0] ), .Z(n18759)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3231_2_lut_rep_577.init = 16'h8888;
    LUT4 i3242_4_lut_3_lut_rep_512_4_lut (.A(n6871[5]), .B(\fcw_r[0] ), 
         .C(n6871[6]), .D(\fcw_r[1] ), .Z(n18694)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3242_4_lut_3_lut_rep_512_4_lut.init = 16'hf880;
    LUT4 i1_2_lut_3_lut (.A(n6871[5]), .B(\fcw_r[0] ), .C(n6871[6]), .Z(n4)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_2_lut_4_lut (.A(\fcw_r[1] ), .B(n18759), .C(n6871[6]), .D(n6871[7]), 
         .Z(n4_adj_839)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_4_lut.init = 16'h17e8;
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count6[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count6[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count6[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count6[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count6[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count6[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count6[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=102, LSE_RLINE=111 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    FD1S3AX fcw_r_ret4_i3 (.D(\fcw_r_15__N_495[8] ), .CK(clk_N_168), .Q(\fcw_r[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret4_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_ret4_i4 (.D(\fcw_r_15__N_495[5] ), .CK(clk_N_168), .Q(fcw_r[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret4_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_ret4_i5 (.D(n16936), .CK(clk_N_168), .Q(fcw_r[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret4_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_ret4_i6 (.D(n15966), .CK(clk_N_168), .Q(n6871[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret4_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_ret4_i7 (.D(n7919[6]), .CK(clk_N_168), .Q(n6871[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret4_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_ret4_i8 (.D(n7920), .CK(clk_N_168), .Q(n6871[7]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret4_i8.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U3
//

module DDS_U3 (\count5[23] , GND_net, \count5[24] , \count_24__N_543[23] , 
            \count_24__N_543[24] , \count5[21] , \count5[22] , \count_24__N_543[21] , 
            \count_24__N_543[22] , \count5[19] , \count5[20] , \count_24__N_543[19] , 
            \count_24__N_543[20] , \count5[17] , \count5[18] , \count_24__N_543[17] , 
            \count_24__N_543[18] , \count5[15] , \count5[16] , \count_24__N_543[15] , 
            \count_24__N_543[16] , \count5[14] , \count_24__N_543[13] , 
            \count_24__N_543[14] , \fcw_r[1] , \count_24__N_543[11] , 
            \count_24__N_543[12] , \count5[1] , clk_N_168, pwm_out2_N_125, 
            n49, n48, n47, n46, n45, n44, n43, n42, n41, n40, 
            n39, n38, n37, n36, n35, n34, n33, n32, n31, n30, 
            n29, n28, n27, n26, \fcw_r[2] , \count_24__N_543[9] , 
            \count_24__N_543[10] , \fcw_r[0] , \count_24__N_543[7] , \count_24__N_543[8] , 
            n18705, n18717, n19839, n8147, n8146, n19840, \count_24__N_543[5] , 
            \count_24__N_543[6] , \count_24__N_543[3] , \count_24__N_543[4] , 
            \count_24__N_543[2] ) /* synthesis syn_module_defined=1 */ ;
    output \count5[23] ;
    input GND_net;
    output \count5[24] ;
    output \count_24__N_543[23] ;
    output \count_24__N_543[24] ;
    output \count5[21] ;
    output \count5[22] ;
    output \count_24__N_543[21] ;
    output \count_24__N_543[22] ;
    output \count5[19] ;
    output \count5[20] ;
    output \count_24__N_543[19] ;
    output \count_24__N_543[20] ;
    output \count5[17] ;
    output \count5[18] ;
    output \count_24__N_543[17] ;
    output \count_24__N_543[18] ;
    output \count5[15] ;
    output \count5[16] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[16] ;
    output \count5[14] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[14] ;
    input \fcw_r[1] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[12] ;
    output \count5[1] ;
    input clk_N_168;
    input pwm_out2_N_125;
    input n49;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    input \fcw_r[2] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[10] ;
    input \fcw_r[0] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[8] ;
    input n18705;
    input n18717;
    input n19839;
    input n8147;
    input n8146;
    input n19840;
    output \count_24__N_543[5] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[3] ;
    output \count_24__N_543[4] ;
    output \count_24__N_543[2] ;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15391, n15390, n15389, n15388, n15387, n15386;
    wire [24:0]count5;   // d:/fpga_project/lattice_diamond/piano/speaker.v(12[33:39])
    
    wire n18723;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    wire [10:0]n6895;
    
    wire n4, n15385, n15384, n18674, n15383, n4_adj_837, n15382, 
        n15381;
    
    CCU2D add_2210_24 (.A0(\count5[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count5[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15391), .S0(\count_24__N_543[23] ), .S1(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_24.INIT0 = 16'h5aaa;
    defparam add_2210_24.INIT1 = 16'h5aaa;
    defparam add_2210_24.INJECT1_0 = "NO";
    defparam add_2210_24.INJECT1_1 = "NO";
    CCU2D add_2210_22 (.A0(\count5[21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count5[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15390), .COUT(n15391), .S0(\count_24__N_543[21] ), 
          .S1(\count_24__N_543[22] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_22.INIT0 = 16'h5aaa;
    defparam add_2210_22.INIT1 = 16'h5aaa;
    defparam add_2210_22.INJECT1_0 = "NO";
    defparam add_2210_22.INJECT1_1 = "NO";
    CCU2D add_2210_20 (.A0(\count5[19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count5[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15389), .COUT(n15390), .S0(\count_24__N_543[19] ), 
          .S1(\count_24__N_543[20] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_20.INIT0 = 16'h5aaa;
    defparam add_2210_20.INIT1 = 16'h5aaa;
    defparam add_2210_20.INJECT1_0 = "NO";
    defparam add_2210_20.INJECT1_1 = "NO";
    CCU2D add_2210_18 (.A0(\count5[17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count5[18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15388), .COUT(n15389), .S0(\count_24__N_543[17] ), 
          .S1(\count_24__N_543[18] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_18.INIT0 = 16'h5aaa;
    defparam add_2210_18.INIT1 = 16'h5aaa;
    defparam add_2210_18.INJECT1_0 = "NO";
    defparam add_2210_18.INJECT1_1 = "NO";
    CCU2D add_2210_16 (.A0(\count5[15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count5[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15387), .COUT(n15388), .S0(\count_24__N_543[15] ), 
          .S1(\count_24__N_543[16] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_16.INIT0 = 16'h5aaa;
    defparam add_2210_16.INIT1 = 16'h5aaa;
    defparam add_2210_16.INJECT1_0 = "NO";
    defparam add_2210_16.INJECT1_1 = "NO";
    CCU2D add_2210_14 (.A0(count5[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count5[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15386), .COUT(n15387), .S0(\count_24__N_543[13] ), .S1(\count_24__N_543[14] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_14.INIT0 = 16'h5aaa;
    defparam add_2210_14.INIT1 = 16'h5aaa;
    defparam add_2210_14.INJECT1_0 = "NO";
    defparam add_2210_14.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(\fcw_r[1] ), .B(n18723), .C(fcw_r[4]), .D(n6895[8]), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_4_lut.init = 16'h17e8;
    CCU2D add_2210_12 (.A0(count5[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count5[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15385), .COUT(n15386), .S0(\count_24__N_543[11] ), .S1(\count_24__N_543[12] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_12.INIT0 = 16'h5aaa;
    defparam add_2210_12.INIT1 = 16'h5aaa;
    defparam add_2210_12.INJECT1_0 = "NO";
    defparam add_2210_12.INJECT1_1 = "NO";
    FD1S3DX count__i1 (.D(n49), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count5[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i1.GSR = "DISABLED";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count5[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count5[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count5[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count5[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count5[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count5[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=91, LSE_RLINE=100 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    CCU2D add_2210_10 (.A0(\fcw_r[2] ), .B0(n4), .C0(count5[9]), .D0(GND_net), 
          .A1(count5[10]), .B1(n18674), .C1(\fcw_r[2] ), .D1(n6895[8]), 
          .CIN(n15384), .COUT(n15385), .S0(\count_24__N_543[9] ), .S1(\count_24__N_543[10] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_10.INIT0 = 16'h9696;
    defparam add_2210_10.INIT1 = 16'h566a;
    defparam add_2210_10.INJECT1_0 = "NO";
    defparam add_2210_10.INJECT1_1 = "NO";
    CCU2D add_2210_8 (.A0(fcw_r[3]), .B0(\fcw_r[0] ), .C0(count5[7]), 
          .D0(GND_net), .A1(\fcw_r[1] ), .B1(n4_adj_837), .C1(count5[8]), 
          .D1(GND_net), .CIN(n15383), .COUT(n15384), .S0(\count_24__N_543[7] ), 
          .S1(\count_24__N_543[8] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_8.INIT0 = 16'h9696;
    defparam add_2210_8.INIT1 = 16'h9696;
    defparam add_2210_8.INJECT1_0 = "NO";
    defparam add_2210_8.INJECT1_1 = "NO";
    FD1S3AX fcw_r_ret6_i2 (.D(n18705), .CK(clk_N_168), .Q(fcw_r[2]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret6_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_ret6_i3 (.D(n18717), .CK(clk_N_168), .Q(fcw_r[3]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret6_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_ret6_i4 (.D(n19839), .CK(clk_N_168), .Q(fcw_r[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret6_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_ret6_i5 (.D(n8147), .CK(clk_N_168), .Q(fcw_r[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret6_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_ret6_i6 (.D(n8146), .CK(clk_N_168), .Q(fcw_r[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret6_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_ret6_i9 (.D(n19840), .CK(clk_N_168), .Q(n6895[8]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret6_i9.GSR = "DISABLED";
    CCU2D add_2210_6 (.A0(count5[5]), .B0(fcw_r[5]), .C0(GND_net), .D0(GND_net), 
          .A1(count5[6]), .B1(fcw_r[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15382), .COUT(n15383), .S0(\count_24__N_543[5] ), .S1(\count_24__N_543[6] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_6.INIT0 = 16'h5666;
    defparam add_2210_6.INIT1 = 16'h5666;
    defparam add_2210_6.INJECT1_0 = "NO";
    defparam add_2210_6.INJECT1_1 = "NO";
    CCU2D add_2210_4 (.A0(count5[3]), .B0(fcw_r[3]), .C0(GND_net), .D0(GND_net), 
          .A1(count5[4]), .B1(fcw_r[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15381), .COUT(n15382), .S0(\count_24__N_543[3] ), .S1(\count_24__N_543[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_4.INIT0 = 16'h5666;
    defparam add_2210_4.INIT1 = 16'h5666;
    defparam add_2210_4.INJECT1_0 = "NO";
    defparam add_2210_4.INJECT1_1 = "NO";
    CCU2D add_2210_2 (.A0(\count5[1] ), .B0(\fcw_r[0] ), .C0(GND_net), 
          .D0(GND_net), .A1(count5[2]), .B1(fcw_r[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15381), .S1(\count_24__N_543[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2210_2.INIT0 = 16'h7000;
    defparam add_2210_2.INIT1 = 16'h5666;
    defparam add_2210_2.INJECT1_0 = "NO";
    defparam add_2210_2.INJECT1_1 = "NO";
    LUT4 i3387_2_lut_rep_541 (.A(fcw_r[3]), .B(\fcw_r[0] ), .Z(n18723)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3387_2_lut_rep_541.init = 16'h8888;
    LUT4 i3398_4_lut_3_lut_rep_492_4_lut (.A(fcw_r[3]), .B(\fcw_r[0] ), 
         .C(fcw_r[4]), .D(\fcw_r[1] ), .Z(n18674)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3398_4_lut_3_lut_rep_492_4_lut.init = 16'hf880;
    LUT4 i1_2_lut_3_lut (.A(fcw_r[3]), .B(\fcw_r[0] ), .C(fcw_r[4]), .Z(n4_adj_837)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    
endmodule
//
// Verilog Description of module DDS_U4
//

module DDS_U4 (\fcw_r[1] , clk_N_168, n18784, \count4[24] , GND_net, 
            n106, \count4[22] , \count4[23] , n108, n107, \count4[20] , 
            \count4[21] , n110, n109, \count4[18] , \count4[19] , 
            n112, n111, \count4[16] , \count4[17] , n114, n113, 
            \count4[14] , \count4[15] , n116, n115, n118, n117, 
            n120, n119, \fcw_r[2] , n122, n121, \fcw_r[0] , n124, 
            n123, n126, n125, n128, n127, n25, n129, pwm_out2_N_125, 
            n132, n18757, \fcw_r_15__N_495[11] , yinjie, n18785, n19846, 
            \yinjie_box[1] , \fcw_r_15__N_527[0] , clk__inv) /* synthesis syn_module_defined=1 */ ;
    output \fcw_r[1] ;
    input clk_N_168;
    input n18784;
    output \count4[24] ;
    input GND_net;
    output n106;
    output \count4[22] ;
    output \count4[23] ;
    output n108;
    output n107;
    output \count4[20] ;
    output \count4[21] ;
    output n110;
    output n109;
    output \count4[18] ;
    output \count4[19] ;
    output n112;
    output n111;
    output \count4[16] ;
    output \count4[17] ;
    output n114;
    output n113;
    output \count4[14] ;
    output \count4[15] ;
    output n116;
    output n115;
    output n118;
    output n117;
    output n120;
    output n119;
    output \fcw_r[2] ;
    output n122;
    output n121;
    input \fcw_r[0] ;
    output n124;
    output n123;
    output n126;
    output n125;
    output n128;
    output n127;
    output n25;
    output n129;
    input pwm_out2_N_125;
    input [24:0]n132;
    input n18757;
    input \fcw_r_15__N_495[11] ;
    input [2:0]yinjie;
    input n18785;
    input n19846;
    input \yinjie_box[1] ;
    input \fcw_r_15__N_527[0] ;
    input clk__inv;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    
    wire n15747, n15746, n15745, n15744, n15743, n15742, n15741;
    wire [24:0]n184;
    
    wire n15740;
    wire [11:0]n6921;
    
    wire n20, n15739, n4, n4_adj_835, n15738;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15737, n15736, n15808;
    wire [9:0]n8293;
    
    wire n8304, n15807, n15806, n18777, n18702;
    
    FD1S3AX fcw_r_ret8_i1 (.D(n18784), .CK(clk_N_168), .Q(\fcw_r[1] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i1.GSR = "DISABLED";
    CCU2D count_2228_add_4_26 (.A0(\count4[24] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15747), .S0(n106));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_26.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_26.INIT1 = 16'h0000;
    defparam count_2228_add_4_26.INJECT1_0 = "NO";
    defparam count_2228_add_4_26.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_24 (.A0(\count4[22] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count4[23] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15746), .COUT(n15747), .S0(n108), .S1(n107));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_24.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_24.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_24.INJECT1_0 = "NO";
    defparam count_2228_add_4_24.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_22 (.A0(\count4[20] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count4[21] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15745), .COUT(n15746), .S0(n110), .S1(n109));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_22.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_22.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_22.INJECT1_0 = "NO";
    defparam count_2228_add_4_22.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_20 (.A0(\count4[18] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count4[19] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15744), .COUT(n15745), .S0(n112), .S1(n111));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_20.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_20.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_20.INJECT1_0 = "NO";
    defparam count_2228_add_4_20.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_18 (.A0(\count4[16] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count4[17] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15743), .COUT(n15744), .S0(n114), .S1(n113));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_18.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_18.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_18.INJECT1_0 = "NO";
    defparam count_2228_add_4_18.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_16 (.A0(\count4[14] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count4[15] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15742), .COUT(n15743), .S0(n116), .S1(n115));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_16.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_16.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_16.INJECT1_0 = "NO";
    defparam count_2228_add_4_16.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_14 (.A0(n184[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n184[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15741), .COUT(n15742), .S0(n118), .S1(n117));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_14.INIT0 = 16'hfaaa;
    defparam count_2228_add_4_14.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_14.INJECT1_0 = "NO";
    defparam count_2228_add_4_14.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_12 (.A0(n6921[10]), .B0(n20), .C0(n184[10]), 
          .D0(GND_net), .A1(n184[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15740), .COUT(n15741), .S0(n120), .S1(n119));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_12.INIT0 = 16'h9696;
    defparam count_2228_add_4_12.INIT1 = 16'hfaaa;
    defparam count_2228_add_4_12.INJECT1_0 = "NO";
    defparam count_2228_add_4_12.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_10 (.A0(\fcw_r[1] ), .B0(n4), .C0(n184[8]), 
          .D0(GND_net), .A1(\fcw_r[2] ), .B1(n4_adj_835), .C1(n184[9]), 
          .D1(GND_net), .CIN(n15739), .COUT(n15740), .S0(n122), .S1(n121));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_10.INIT0 = 16'h9696;
    defparam count_2228_add_4_10.INIT1 = 16'h9696;
    defparam count_2228_add_4_10.INJECT1_0 = "NO";
    defparam count_2228_add_4_10.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_8 (.A0(fcw_r[6]), .B0(n184[6]), .C0(GND_net), 
          .D0(GND_net), .A1(n6921[7]), .B1(\fcw_r[0] ), .C1(n184[7]), 
          .D1(GND_net), .CIN(n15738), .COUT(n15739), .S0(n124), .S1(n123));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_8.INIT0 = 16'h5666;
    defparam count_2228_add_4_8.INIT1 = 16'h9696;
    defparam count_2228_add_4_8.INJECT1_0 = "NO";
    defparam count_2228_add_4_8.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_6 (.A0(fcw_r[4]), .B0(n184[4]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[5]), .B1(n184[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15737), .COUT(n15738), .S0(n126), .S1(n125));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_6.INIT0 = 16'h5666;
    defparam count_2228_add_4_6.INIT1 = 16'h5666;
    defparam count_2228_add_4_6.INJECT1_0 = "NO";
    defparam count_2228_add_4_6.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_4 (.A0(\fcw_r[2] ), .B0(n184[2]), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[0] ), .B1(n184[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15736), .COUT(n15737), .S0(n128), .S1(n127));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_4.INIT0 = 16'h5666;
    defparam count_2228_add_4_4.INIT1 = 16'h5666;
    defparam count_2228_add_4_4.INJECT1_0 = "NO";
    defparam count_2228_add_4_4.INJECT1_1 = "NO";
    CCU2D count_2228_add_4_2 (.A0(\fcw_r[0] ), .B0(n25), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[1] ), .B1(n184[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15736), .S1(n129));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228_add_4_2.INIT0 = 16'h7000;
    defparam count_2228_add_4_2.INIT1 = 16'h5666;
    defparam count_2228_add_4_2.INJECT1_0 = "NO";
    defparam count_2228_add_4_2.INJECT1_1 = "NO";
    FD1S3DX count_2228__i0 (.D(n132[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n25)) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i0.GSR = "DISABLED";
    CCU2D add_3609_7 (.A0(n18757), .B0(\fcw_r_15__N_495[11] ), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15808), .S0(n8293[9]), .S1(n8304));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3609_7.INIT0 = 16'h7888;
    defparam add_3609_7.INIT1 = 16'h0000;
    defparam add_3609_7.INJECT1_0 = "NO";
    defparam add_3609_7.INJECT1_1 = "NO";
    CCU2D add_3609_5 (.A0(yinjie[2]), .B0(n18785), .C0(n18784), .D0(n19846), 
          .A1(n18757), .B1(\fcw_r_15__N_495[11] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15807), .COUT(n15808), .S0(n8293[7]), .S1(n8293[8]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3609_5.INIT0 = 16'hf078;
    defparam add_3609_5.INIT1 = 16'h9666;
    defparam add_3609_5.INJECT1_0 = "NO";
    defparam add_3609_5.INJECT1_1 = "NO";
    CCU2D add_3609_3 (.A0(yinjie[2]), .B0(n19846), .C0(\yinjie_box[1] ), 
          .D0(yinjie[1]), .A1(yinjie[2]), .B1(yinjie[0]), .C1(\fcw_r_15__N_527[0] ), 
          .D1(n19846), .CIN(n15806), .COUT(n15807), .S0(n8293[5]), .S1(n8293[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3609_3.INIT0 = 16'hd1e2;
    defparam add_3609_3.INIT1 = 16'hf066;
    defparam add_3609_3.INJECT1_0 = "NO";
    defparam add_3609_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(\fcw_r[1] ), .B(n18777), .C(n6921[8]), .D(n6921[9]), 
         .Z(n4_adj_835)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_4_lut.init = 16'h17e8;
    CCU2D add_3609_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n18784), .B1(n19846), .C1(\fcw_r_15__N_527[0] ), .D1(yinjie[0]), 
          .COUT(n15806), .S1(n8293[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3609_1.INIT0 = 16'hF000;
    defparam add_3609_1.INIT1 = 16'h596a;
    defparam add_3609_1.INJECT1_0 = "NO";
    defparam add_3609_1.INJECT1_1 = "NO";
    LUT4 i3521_2_lut_rep_595 (.A(n6921[7]), .B(\fcw_r[0] ), .Z(n18777)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3521_2_lut_rep_595.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(n6921[7]), .B(\fcw_r[0] ), .C(n6921[8]), .Z(n4)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 i3532_4_lut_3_lut_rep_520_4_lut (.A(n6921[7]), .B(\fcw_r[0] ), 
         .C(n6921[8]), .D(\fcw_r[1] ), .Z(n18702)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3532_4_lut_3_lut_rep_520_4_lut.init = 16'hf880;
    FD1S3AX fcw_r_ret8_i2 (.D(n18757), .CK(clk_N_168), .Q(\fcw_r[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i4 (.D(n8293[4]), .CK(clk_N_168), .Q(fcw_r[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i5 (.D(n8293[5]), .CK(clk_N_168), .Q(fcw_r[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i6 (.D(n8293[6]), .CK(clk_N_168), .Q(fcw_r[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i7 (.D(n8293[7]), .CK(clk_N_168), .Q(n6921[7]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i8 (.D(n8293[8]), .CK(clk_N_168), .Q(n6921[8]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i8.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i9 (.D(n8293[9]), .CK(clk_N_168), .Q(n6921[9]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i9.GSR = "DISABLED";
    FD1S3AX fcw_r_ret8_i10 (.D(n8304), .CK(clk_N_168), .Q(n6921[10]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret8_i10.GSR = "DISABLED";
    FD1S3DX count_2228__i1 (.D(n132[1]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i1.GSR = "DISABLED";
    FD1S3DX count_2228__i2 (.D(n132[2]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i2.GSR = "DISABLED";
    FD1S3DX count_2228__i3 (.D(n132[3]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i3.GSR = "DISABLED";
    FD1S3DX count_2228__i4 (.D(n132[4]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i4.GSR = "DISABLED";
    FD1S3DX count_2228__i5 (.D(n132[5]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i5.GSR = "DISABLED";
    FD1S3DX count_2228__i6 (.D(n132[6]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i6.GSR = "DISABLED";
    FD1S3DX count_2228__i7 (.D(n132[7]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i7.GSR = "DISABLED";
    FD1S3DX count_2228__i8 (.D(n132[8]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i8.GSR = "DISABLED";
    FD1S3DX count_2228__i9 (.D(n132[9]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i9.GSR = "DISABLED";
    FD1S3DX count_2228__i10 (.D(n132[10]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i10.GSR = "DISABLED";
    FD1S3DX count_2228__i11 (.D(n132[11]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i11.GSR = "DISABLED";
    FD1S3DX count_2228__i12 (.D(n132[12]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i12.GSR = "DISABLED";
    FD1S3DX count_2228__i13 (.D(n132[13]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i13.GSR = "DISABLED";
    FD1S3DX count_2228__i14 (.D(n132[14]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[14] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i14.GSR = "DISABLED";
    FD1S3DX count_2228__i15 (.D(n132[15]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[15] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i15.GSR = "DISABLED";
    FD1S3DX count_2228__i16 (.D(n132[16]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[16] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i16.GSR = "DISABLED";
    FD1S3DX count_2228__i17 (.D(n132[17]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[17] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i17.GSR = "DISABLED";
    FD1S3DX count_2228__i18 (.D(n132[18]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[18] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i18.GSR = "DISABLED";
    FD1S3DX count_2228__i19 (.D(n132[19]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[19] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i19.GSR = "DISABLED";
    FD1S3DX count_2228__i20 (.D(n132[20]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[20] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i20.GSR = "DISABLED";
    FD1S3DX count_2228__i21 (.D(n132[21]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[21] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i21.GSR = "DISABLED";
    FD1S3DX count_2228__i22 (.D(n132[22]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[22] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i22.GSR = "DISABLED";
    FD1S3DX count_2228__i23 (.D(n132[23]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[23] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i23.GSR = "DISABLED";
    FD1S3DX count_2228__i24 (.D(n132[24]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count4[24] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2228__i24.GSR = "DISABLED";
    LUT4 i3539_4_lut_3_lut (.A(\fcw_r[2] ), .B(n18702), .C(n6921[9]), 
         .Z(n20)) /* synthesis lut_function=(A (B+(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3539_4_lut_3_lut.init = 16'he8e8;
    
endmodule
//
// Verilog Description of module DDS_U5
//

module DDS_U5 (\fcw_r[0] , clk_N_168, n18785, \count3[24] , GND_net, 
            n106, \count3[22] , \count3[23] , n108, n107, \count3[20] , 
            \count3[21] , n110, n109, \count3[18] , \count3[19] , 
            n112, n111, \count3[16] , \count3[17] , n114, n113, 
            \count3[14] , \count3[15] , n116, n115, n118, n117, 
            \fcw_r[2] , n120, n119, \fcw_r[1] , n122, n121, n124, 
            n123, n126, n125, \fcw_r[4] , n128, n127, n25, n129, 
            pwm_out2_N_125, n132, \yinjie[2] , n19846, n18784, \fcw_r_15__N_495[11] , 
            \fcw_r_15__N_495[9] , \fcw_r_15__N_527[0] , \yinjie[0] , clk__inv) /* synthesis syn_module_defined=1 */ ;
    output \fcw_r[0] ;
    input clk_N_168;
    input n18785;
    output \count3[24] ;
    input GND_net;
    output n106;
    output \count3[22] ;
    output \count3[23] ;
    output n108;
    output n107;
    output \count3[20] ;
    output \count3[21] ;
    output n110;
    output n109;
    output \count3[18] ;
    output \count3[19] ;
    output n112;
    output n111;
    output \count3[16] ;
    output \count3[17] ;
    output n114;
    output n113;
    output \count3[14] ;
    output \count3[15] ;
    output n116;
    output n115;
    output n118;
    output n117;
    input \fcw_r[2] ;
    output n120;
    output n119;
    input \fcw_r[1] ;
    output n122;
    output n121;
    output n124;
    output n123;
    output n126;
    output n125;
    input \fcw_r[4] ;
    output n128;
    output n127;
    output n25;
    output n129;
    input pwm_out2_N_125;
    input [24:0]n132;
    input \yinjie[2] ;
    input n19846;
    input n18784;
    input \fcw_r_15__N_495[11] ;
    input \fcw_r_15__N_495[9] ;
    input \fcw_r_15__N_527[0] ;
    input \yinjie[0] ;
    input clk__inv;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    
    wire n15760, n15759, n15758, n15757, n15756, n15755, n15754;
    wire [24:0]n184;
    
    wire n15753, n18703;
    wire [11:0]n6843;
    
    wire n15752, n4, n4_adj_833, n15751;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15750, n15749, n15498;
    wire [8:0]n8382;
    
    wire n8392, n15497, n15496, n18778;
    
    FD1S3AX fcw_r_ret2_i1 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[0] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i1.GSR = "DISABLED";
    CCU2D count_2227_add_4_26 (.A0(\count3[24] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15760), .S0(n106));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_26.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_26.INIT1 = 16'h0000;
    defparam count_2227_add_4_26.INJECT1_0 = "NO";
    defparam count_2227_add_4_26.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_24 (.A0(\count3[22] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count3[23] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15759), .COUT(n15760), .S0(n108), .S1(n107));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_24.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_24.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_24.INJECT1_0 = "NO";
    defparam count_2227_add_4_24.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_22 (.A0(\count3[20] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count3[21] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15758), .COUT(n15759), .S0(n110), .S1(n109));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_22.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_22.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_22.INJECT1_0 = "NO";
    defparam count_2227_add_4_22.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_20 (.A0(\count3[18] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count3[19] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15757), .COUT(n15758), .S0(n112), .S1(n111));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_20.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_20.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_20.INJECT1_0 = "NO";
    defparam count_2227_add_4_20.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_18 (.A0(\count3[16] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count3[17] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15756), .COUT(n15757), .S0(n114), .S1(n113));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_18.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_18.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_18.INJECT1_0 = "NO";
    defparam count_2227_add_4_18.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_16 (.A0(\count3[14] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count3[15] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15755), .COUT(n15756), .S0(n116), .S1(n115));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_16.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_16.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_16.INJECT1_0 = "NO";
    defparam count_2227_add_4_16.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_14 (.A0(n184[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n184[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15754), .COUT(n15755), .S0(n118), .S1(n117));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_14.INIT0 = 16'hfaaa;
    defparam count_2227_add_4_14.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_14.INJECT1_0 = "NO";
    defparam count_2227_add_4_14.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_12 (.A0(n184[10]), .B0(n18703), .C0(\fcw_r[2] ), 
          .D0(n6843[9]), .A1(n184[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15753), .COUT(n15754), .S0(n120), .S1(n119));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_12.INIT0 = 16'h566a;
    defparam count_2227_add_4_12.INIT1 = 16'hfaaa;
    defparam count_2227_add_4_12.INJECT1_0 = "NO";
    defparam count_2227_add_4_12.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_10 (.A0(\fcw_r[1] ), .B0(n4), .C0(n184[8]), 
          .D0(GND_net), .A1(\fcw_r[2] ), .B1(n4_adj_833), .C1(n184[9]), 
          .D1(GND_net), .CIN(n15752), .COUT(n15753), .S0(n122), .S1(n121));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_10.INIT0 = 16'h9696;
    defparam count_2227_add_4_10.INIT1 = 16'h9696;
    defparam count_2227_add_4_10.INJECT1_0 = "NO";
    defparam count_2227_add_4_10.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_8 (.A0(fcw_r[6]), .B0(n184[6]), .C0(GND_net), 
          .D0(GND_net), .A1(n6843[7]), .B1(\fcw_r[0] ), .C1(n184[7]), 
          .D1(GND_net), .CIN(n15751), .COUT(n15752), .S0(n124), .S1(n123));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_8.INIT0 = 16'h5666;
    defparam count_2227_add_4_8.INIT1 = 16'h9696;
    defparam count_2227_add_4_8.INJECT1_0 = "NO";
    defparam count_2227_add_4_8.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_6 (.A0(fcw_r[4]), .B0(n184[4]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[5]), .B1(n184[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15750), .COUT(n15751), .S0(n126), .S1(n125));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_6.INIT0 = 16'h5666;
    defparam count_2227_add_4_6.INIT1 = 16'h5666;
    defparam count_2227_add_4_6.INJECT1_0 = "NO";
    defparam count_2227_add_4_6.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_4 (.A0(\fcw_r[4] ), .B0(n184[2]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[3]), .B1(n184[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15749), .COUT(n15750), .S0(n128), .S1(n127));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_4.INIT0 = 16'h5666;
    defparam count_2227_add_4_4.INIT1 = 16'h5666;
    defparam count_2227_add_4_4.INJECT1_0 = "NO";
    defparam count_2227_add_4_4.INJECT1_1 = "NO";
    CCU2D count_2227_add_4_2 (.A0(\fcw_r[0] ), .B0(n25), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[1] ), .B1(n184[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15749), .S1(n129));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227_add_4_2.INIT0 = 16'h7000;
    defparam count_2227_add_4_2.INIT1 = 16'h5666;
    defparam count_2227_add_4_2.INJECT1_0 = "NO";
    defparam count_2227_add_4_2.INJECT1_1 = "NO";
    FD1S3DX count_2227__i0 (.D(n132[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n25)) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i0.GSR = "DISABLED";
    CCU2D add_3687_7 (.A0(\yinjie[2] ), .B0(n19846), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15498), 
          .S0(n8382[8]), .S1(n8392));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3687_7.INIT0 = 16'hd222;
    defparam add_3687_7.INIT1 = 16'h0000;
    defparam add_3687_7.INJECT1_0 = "NO";
    defparam add_3687_7.INJECT1_1 = "NO";
    CCU2D add_3687_5 (.A0(n18785), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n18784), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15497), 
          .COUT(n15498), .S0(n8382[6]), .S1(n8382[7]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3687_5.INIT0 = 16'hfaaa;
    defparam add_3687_5.INIT1 = 16'hfaaa;
    defparam add_3687_5.INJECT1_0 = "NO";
    defparam add_3687_5.INJECT1_1 = "NO";
    CCU2D add_3687_3 (.A0(n18784), .B0(\yinjie[2] ), .C0(\fcw_r_15__N_495[11] ), 
          .D0(n19846), .A1(\yinjie[2] ), .B1(n19846), .C1(\fcw_r_15__N_495[11] ), 
          .D1(GND_net), .CIN(n15496), .COUT(n15497), .S0(n8382[4]), 
          .S1(n8382[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3687_3.INIT0 = 16'h5a96;
    defparam add_3687_3.INIT1 = 16'hd2d2;
    defparam add_3687_3.INJECT1_0 = "NO";
    defparam add_3687_3.INJECT1_1 = "NO";
    CCU2D add_3687_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\fcw_r_15__N_495[9] ), .B1(n19846), .C1(\fcw_r_15__N_527[0] ), 
          .D1(\yinjie[0] ), .COUT(n15496), .S1(n8382[3]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3687_1.INIT0 = 16'hF000;
    defparam add_3687_1.INIT1 = 16'h596a;
    defparam add_3687_1.INJECT1_0 = "NO";
    defparam add_3687_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(\fcw_r[1] ), .B(n18778), .C(n6843[8]), .D(n6843[9]), 
         .Z(n4_adj_833)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_4_lut.init = 16'h17e8;
    LUT4 i3662_2_lut_rep_596 (.A(n6843[7]), .B(\fcw_r[0] ), .Z(n18778)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3662_2_lut_rep_596.init = 16'h8888;
    LUT4 i3673_4_lut_3_lut_rep_521_4_lut (.A(n6843[7]), .B(\fcw_r[0] ), 
         .C(n6843[8]), .D(\fcw_r[1] ), .Z(n18703)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3673_4_lut_3_lut_rep_521_4_lut.init = 16'hf880;
    LUT4 i1_2_lut_3_lut (.A(n6843[7]), .B(\fcw_r[0] ), .C(n6843[8]), .Z(n4)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    FD1S3AX fcw_r_ret2_i4 (.D(n8382[3]), .CK(clk_N_168), .Q(fcw_r[3]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_ret2_i5 (.D(n8382[4]), .CK(clk_N_168), .Q(fcw_r[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_ret2_i6 (.D(n8382[5]), .CK(clk_N_168), .Q(fcw_r[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_ret2_i7 (.D(n8382[6]), .CK(clk_N_168), .Q(fcw_r[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_ret2_i8 (.D(n8382[7]), .CK(clk_N_168), .Q(n6843[7]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i8.GSR = "DISABLED";
    FD1S3AX fcw_r_ret2_i9 (.D(n8382[8]), .CK(clk_N_168), .Q(n6843[8]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i9.GSR = "DISABLED";
    FD1S3AX fcw_r_ret2_i10 (.D(n8392), .CK(clk_N_168), .Q(n6843[9]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret2_i10.GSR = "DISABLED";
    FD1S3DX count_2227__i1 (.D(n132[1]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i1.GSR = "DISABLED";
    FD1S3DX count_2227__i2 (.D(n132[2]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i2.GSR = "DISABLED";
    FD1S3DX count_2227__i3 (.D(n132[3]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i3.GSR = "DISABLED";
    FD1S3DX count_2227__i4 (.D(n132[4]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i4.GSR = "DISABLED";
    FD1S3DX count_2227__i5 (.D(n132[5]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i5.GSR = "DISABLED";
    FD1S3DX count_2227__i6 (.D(n132[6]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i6.GSR = "DISABLED";
    FD1S3DX count_2227__i7 (.D(n132[7]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i7.GSR = "DISABLED";
    FD1S3DX count_2227__i8 (.D(n132[8]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i8.GSR = "DISABLED";
    FD1S3DX count_2227__i9 (.D(n132[9]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i9.GSR = "DISABLED";
    FD1S3DX count_2227__i10 (.D(n132[10]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i10.GSR = "DISABLED";
    FD1S3DX count_2227__i11 (.D(n132[11]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i11.GSR = "DISABLED";
    FD1S3DX count_2227__i12 (.D(n132[12]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i12.GSR = "DISABLED";
    FD1S3DX count_2227__i13 (.D(n132[13]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i13.GSR = "DISABLED";
    FD1S3DX count_2227__i14 (.D(n132[14]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[14] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i14.GSR = "DISABLED";
    FD1S3DX count_2227__i15 (.D(n132[15]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[15] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i15.GSR = "DISABLED";
    FD1S3DX count_2227__i16 (.D(n132[16]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[16] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i16.GSR = "DISABLED";
    FD1S3DX count_2227__i17 (.D(n132[17]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[17] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i17.GSR = "DISABLED";
    FD1S3DX count_2227__i18 (.D(n132[18]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[18] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i18.GSR = "DISABLED";
    FD1S3DX count_2227__i19 (.D(n132[19]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[19] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i19.GSR = "DISABLED";
    FD1S3DX count_2227__i20 (.D(n132[20]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[20] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i20.GSR = "DISABLED";
    FD1S3DX count_2227__i21 (.D(n132[21]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[21] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i21.GSR = "DISABLED";
    FD1S3DX count_2227__i22 (.D(n132[22]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[22] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i22.GSR = "DISABLED";
    FD1S3DX count_2227__i23 (.D(n132[23]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[23] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i23.GSR = "DISABLED";
    FD1S3DX count_2227__i24 (.D(n132[24]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count3[24] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2227__i24.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U6
//

module DDS_U6 (clk_N_168, n18784, \count2[23] , GND_net, \count2[24] , 
            \count_24__N_543[23] , \count_24__N_543[24] , \yinjie[1] , 
            n19846, \yinjie[2] , n19840, \count2[21] , \count2[22] , 
            \count_24__N_543[21] , \count_24__N_543[22] , \count2[19] , 
            \count2[20] , \count_24__N_543[19] , \count_24__N_543[20] , 
            \count2[17] , \count2[18] , \count_24__N_543[17] , \count_24__N_543[18] , 
            \count2[15] , \count2[16] , \count_24__N_543[15] , \count_24__N_543[16] , 
            \count2[14] , \count_24__N_543[13] , \count_24__N_543[14] , 
            \count_24__N_543[11] , \count_24__N_543[12] , \count_24__N_543[9] , 
            \count_24__N_543[10] , \count_24__N_543[7] , \count_24__N_543[8] , 
            n18757, \fcw_r[6] , n18785, n18705, n18717, n19839, 
            \yinjie_box[1] , n18716, \count2[1] , pwm_out2_N_125, n49, 
            n48, n47, n46, n45, n44, n43, n42, n41, n40, n39, 
            n38, n37, n36, n35, n34, n33, n32, n31, n30, n29, 
            n28, n27, n26, \count_24__N_543[5] , \count_24__N_543[6] , 
            \count_24__N_543[3] , \count_24__N_543[4] , \count_24__N_543[2] , 
            n18608, n7920) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output n18784;
    output \count2[23] ;
    input GND_net;
    output \count2[24] ;
    output \count_24__N_543[23] ;
    output \count_24__N_543[24] ;
    input \yinjie[1] ;
    input n19846;
    input \yinjie[2] ;
    output n19840;
    output \count2[21] ;
    output \count2[22] ;
    output \count_24__N_543[21] ;
    output \count_24__N_543[22] ;
    output \count2[19] ;
    output \count2[20] ;
    output \count_24__N_543[19] ;
    output \count_24__N_543[20] ;
    output \count2[17] ;
    output \count2[18] ;
    output \count_24__N_543[17] ;
    output \count_24__N_543[18] ;
    output \count2[15] ;
    output \count2[16] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[16] ;
    output \count2[14] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[14] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[12] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[10] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[8] ;
    input n18757;
    output \fcw_r[6] ;
    input n18785;
    output n18705;
    input n18717;
    input n19839;
    input \yinjie_box[1] ;
    output n18716;
    output \count2[1] ;
    input pwm_out2_N_125;
    input n49;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    output \count_24__N_543[5] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[3] ;
    output \count_24__N_543[4] ;
    output \count_24__N_543[2] ;
    input n18608;
    output n7920;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15494, n15493, n15492, n15491, n15490, n15489;
    wire [24:0]count2;   // d:/fpga_project/lattice_diamond/piano/speaker.v(11[34:40])
    
    wire n15488, n15487, n15486, n15485, n15484;
    
    FD1S3AX fcw_r_i1 (.D(n18784), .CK(clk_N_168), .Q(fcw_r[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D add_2209_24 (.A0(\count2[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count2[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15494), .S0(\count_24__N_543[23] ), .S1(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_24.INIT0 = 16'h5aaa;
    defparam add_2209_24.INIT1 = 16'h5aaa;
    defparam add_2209_24.INJECT1_0 = "NO";
    defparam add_2209_24.INJECT1_1 = "NO";
    LUT4 i4027_3_lut_4_lut_3_lut (.A(\yinjie[1] ), .B(n19846), .C(\yinjie[2] ), 
         .Z(n19840)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i4027_3_lut_4_lut_3_lut.init = 16'h2020;
    CCU2D add_2209_22 (.A0(\count2[21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count2[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15493), .COUT(n15494), .S0(\count_24__N_543[21] ), 
          .S1(\count_24__N_543[22] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_22.INIT0 = 16'h5aaa;
    defparam add_2209_22.INIT1 = 16'h5aaa;
    defparam add_2209_22.INJECT1_0 = "NO";
    defparam add_2209_22.INJECT1_1 = "NO";
    CCU2D add_2209_20 (.A0(\count2[19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count2[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15492), .COUT(n15493), .S0(\count_24__N_543[19] ), 
          .S1(\count_24__N_543[20] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_20.INIT0 = 16'h5aaa;
    defparam add_2209_20.INIT1 = 16'h5aaa;
    defparam add_2209_20.INJECT1_0 = "NO";
    defparam add_2209_20.INJECT1_1 = "NO";
    CCU2D add_2209_18 (.A0(\count2[17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count2[18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15491), .COUT(n15492), .S0(\count_24__N_543[17] ), 
          .S1(\count_24__N_543[18] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_18.INIT0 = 16'h5aaa;
    defparam add_2209_18.INIT1 = 16'h5aaa;
    defparam add_2209_18.INJECT1_0 = "NO";
    defparam add_2209_18.INJECT1_1 = "NO";
    CCU2D add_2209_16 (.A0(\count2[15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count2[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15490), .COUT(n15491), .S0(\count_24__N_543[15] ), 
          .S1(\count_24__N_543[16] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_16.INIT0 = 16'h5aaa;
    defparam add_2209_16.INIT1 = 16'h5aaa;
    defparam add_2209_16.INJECT1_0 = "NO";
    defparam add_2209_16.INJECT1_1 = "NO";
    CCU2D add_2209_14 (.A0(count2[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count2[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15489), .COUT(n15490), .S0(\count_24__N_543[13] ), .S1(\count_24__N_543[14] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_14.INIT0 = 16'h5aaa;
    defparam add_2209_14.INIT1 = 16'h5aaa;
    defparam add_2209_14.INJECT1_0 = "NO";
    defparam add_2209_14.INJECT1_1 = "NO";
    CCU2D add_2209_12 (.A0(count2[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count2[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15488), .COUT(n15489), .S0(\count_24__N_543[11] ), .S1(\count_24__N_543[12] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_12.INIT0 = 16'h5aaa;
    defparam add_2209_12.INIT1 = 16'h5aaa;
    defparam add_2209_12.INJECT1_0 = "NO";
    defparam add_2209_12.INJECT1_1 = "NO";
    CCU2D add_2209_10 (.A0(count2[9]), .B0(fcw_r[9]), .C0(GND_net), .D0(GND_net), 
          .A1(count2[10]), .B1(fcw_r[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15487), .COUT(n15488), .S0(\count_24__N_543[9] ), .S1(\count_24__N_543[10] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_10.INIT0 = 16'h5666;
    defparam add_2209_10.INIT1 = 16'h5666;
    defparam add_2209_10.INJECT1_0 = "NO";
    defparam add_2209_10.INJECT1_1 = "NO";
    CCU2D add_2209_8 (.A0(count2[7]), .B0(fcw_r[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count2[8]), .B1(fcw_r[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15486), .COUT(n15487), .S0(\count_24__N_543[7] ), .S1(\count_24__N_543[8] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_8.INIT0 = 16'h5666;
    defparam add_2209_8.INIT1 = 16'h5666;
    defparam add_2209_8.INJECT1_0 = "NO";
    defparam add_2209_8.INJECT1_1 = "NO";
    FD1S3AX fcw_r_i2 (.D(n18757), .CK(clk_N_168), .Q(fcw_r[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_i4 (.D(n18705), .CK(clk_N_168), .Q(fcw_r[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_i5 (.D(n18717), .CK(clk_N_168), .Q(fcw_r[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_i6 (.D(n19839), .CK(clk_N_168), .Q(fcw_r[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_i7 (.D(n19840), .CK(clk_N_168), .Q(fcw_r[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i7.GSR = "DISABLED";
    LUT4 mux_2173_i2_3_lut_rep_602 (.A(\yinjie[1] ), .B(\yinjie_box[1] ), 
         .C(n19846), .Z(n18784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam mux_2173_i2_3_lut_rep_602.init = 16'hcaca;
    LUT4 i3448_2_lut_rep_523_4_lut (.A(\yinjie[1] ), .B(\yinjie_box[1] ), 
         .C(n19846), .D(n18785), .Z(n18705)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3448_2_lut_rep_523_4_lut.init = 16'h35ca;
    LUT4 i10328_2_lut_rep_534_4_lut (.A(\yinjie[1] ), .B(\yinjie_box[1] ), 
         .C(n19846), .D(n18785), .Z(n18716)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i10328_2_lut_rep_534_4_lut.init = 16'h00ca;
    FD1S3DX count__i1 (.D(n49), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count2[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i1.GSR = "DISABLED";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count2[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count2[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count2[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count2[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count2[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count2[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=58, LSE_RLINE=67 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    CCU2D add_2209_6 (.A0(count2[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count2[6]), .B1(\fcw_r[6] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15485), .COUT(n15486), .S0(\count_24__N_543[5] ), .S1(\count_24__N_543[6] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_6.INIT0 = 16'h5aaa;
    defparam add_2209_6.INIT1 = 16'h5666;
    defparam add_2209_6.INJECT1_0 = "NO";
    defparam add_2209_6.INJECT1_1 = "NO";
    CCU2D add_2209_4 (.A0(count2[3]), .B0(fcw_r[3]), .C0(GND_net), .D0(GND_net), 
          .A1(count2[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15484), .COUT(n15485), .S0(\count_24__N_543[3] ), .S1(\count_24__N_543[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_4.INIT0 = 16'h5666;
    defparam add_2209_4.INIT1 = 16'h5aaa;
    defparam add_2209_4.INJECT1_0 = "NO";
    defparam add_2209_4.INJECT1_1 = "NO";
    CCU2D add_2209_2 (.A0(\count2[1] ), .B0(\fcw_r[6] ), .C0(GND_net), 
          .D0(GND_net), .A1(count2[2]), .B1(fcw_r[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15484), .S1(\count_24__N_543[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2209_2.INIT0 = 16'h7000;
    defparam add_2209_2.INIT1 = 16'h5666;
    defparam add_2209_2.INJECT1_0 = "NO";
    defparam add_2209_2.INJECT1_1 = "NO";
    LUT4 i4155_3_lut_4_lut_4_lut (.A(n18757), .B(n18784), .C(n18785), 
         .D(n18608), .Z(n7920)) /* synthesis lut_function=(A (B+(D))+!A (B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i4155_3_lut_4_lut_4_lut.init = 16'hea88;
    
endmodule
//
// Verilog Description of module DDS_U7
//

module DDS_U7 (n19846, \fcw_r[0] , clk_N_168, n18785, \count1[24] , 
            GND_net, n106, \count1[22] , \count1[23] , n108, n107, 
            \count1[20] , \count1[21] , n110, n109, \count1[18] , 
            \count1[19] , n112, n111, \count1[16] , \count1[17] , 
            n114, n113, \count1[14] , \count1[15] , n116, n115, 
            n118, n117, \fcw_r[10] , n120, n119, \fcw_r[8] , \fcw_r[9] , 
            n122, n121, \fcw_r[6] , \fcw_r[7] , n124, n123, \fcw_r[4] , 
            \fcw_r[5] , n126, n125, \fcw_r[2] , \fcw_r[3] , n128, 
            n127, n25, \fcw_r[1] , n129, yinjie, \yinjie_box[1] , 
            \fcw_r_15__N_527[0] , pwm_out2_N_125, n132, stat, \fcw_r_15__N_495[8] , 
            clk__inv) /* synthesis syn_module_defined=1 */ ;
    input n19846;
    output \fcw_r[0] ;
    input clk_N_168;
    output n18785;
    output \count1[24] ;
    input GND_net;
    output n106;
    output \count1[22] ;
    output \count1[23] ;
    output n108;
    output n107;
    output \count1[20] ;
    output \count1[21] ;
    output n110;
    output n109;
    output \count1[18] ;
    output \count1[19] ;
    output n112;
    output n111;
    output \count1[16] ;
    output \count1[17] ;
    output n114;
    output n113;
    output \count1[14] ;
    output \count1[15] ;
    output n116;
    output n115;
    output n118;
    output n117;
    output \fcw_r[10] ;
    output n120;
    output n119;
    output \fcw_r[8] ;
    output \fcw_r[9] ;
    output n122;
    output n121;
    output \fcw_r[6] ;
    output \fcw_r[7] ;
    output n124;
    output n123;
    output \fcw_r[4] ;
    output \fcw_r[5] ;
    output n126;
    output n125;
    output \fcw_r[2] ;
    output \fcw_r[3] ;
    output n128;
    output n127;
    output n25;
    output \fcw_r[1] ;
    output n129;
    input [2:0]yinjie;
    input \yinjie_box[1] ;
    input \fcw_r_15__N_527[0] ;
    input pwm_out2_N_125;
    input [24:0]n132;
    input stat;
    output \fcw_r_15__N_495[8] ;
    input clk__inv;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire [9:0]n7610;
    wire [18:0]fcw_r_15__N_527;
    wire [15:0]fcw_r_15__N_495;
    
    wire n15773, n15772, n15771, n15770, n15769, n15768, n15767;
    wire [24:0]n184;
    
    wire n15766, n15765, n15764, n15763, n15762, n15512, n7621, 
        n15511, n15510, n8, n15509, n9471;
    wire [10:0]n7597;
    
    wire n18861, n18860, n15802, n15801, n15800;
    
    PFUMX mux_1493_i2 (.BLUT(n7610[1]), .ALUT(fcw_r_15__N_527[1]), .C0(n19846), 
          .Z(fcw_r_15__N_495[1]));
    FD1S3AX fcw_r_i1 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D count_2226_add_4_26 (.A0(\count1[24] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15773), .S0(n106));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_26.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_26.INIT1 = 16'h0000;
    defparam count_2226_add_4_26.INJECT1_0 = "NO";
    defparam count_2226_add_4_26.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_24 (.A0(\count1[22] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count1[23] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15772), .COUT(n15773), .S0(n108), .S1(n107));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_24.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_24.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_24.INJECT1_0 = "NO";
    defparam count_2226_add_4_24.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_22 (.A0(\count1[20] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count1[21] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15771), .COUT(n15772), .S0(n110), .S1(n109));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_22.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_22.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_22.INJECT1_0 = "NO";
    defparam count_2226_add_4_22.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_20 (.A0(\count1[18] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count1[19] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15770), .COUT(n15771), .S0(n112), .S1(n111));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_20.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_20.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_20.INJECT1_0 = "NO";
    defparam count_2226_add_4_20.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_18 (.A0(\count1[16] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count1[17] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15769), .COUT(n15770), .S0(n114), .S1(n113));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_18.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_18.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_18.INJECT1_0 = "NO";
    defparam count_2226_add_4_18.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_16 (.A0(\count1[14] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count1[15] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15768), .COUT(n15769), .S0(n116), .S1(n115));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_16.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_16.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_16.INJECT1_0 = "NO";
    defparam count_2226_add_4_16.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_14 (.A0(n184[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n184[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15767), .COUT(n15768), .S0(n118), .S1(n117));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_14.INIT0 = 16'hfaaa;
    defparam count_2226_add_4_14.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_14.INJECT1_0 = "NO";
    defparam count_2226_add_4_14.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_12 (.A0(\fcw_r[10] ), .B0(n184[10]), .C0(GND_net), 
          .D0(GND_net), .A1(n184[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15766), .COUT(n15767), .S0(n120), .S1(n119));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_12.INIT0 = 16'h5666;
    defparam count_2226_add_4_12.INIT1 = 16'hfaaa;
    defparam count_2226_add_4_12.INJECT1_0 = "NO";
    defparam count_2226_add_4_12.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_10 (.A0(\fcw_r[8] ), .B0(n184[8]), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[9] ), .B1(n184[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15765), .COUT(n15766), .S0(n122), .S1(n121));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_10.INIT0 = 16'h5666;
    defparam count_2226_add_4_10.INIT1 = 16'h5666;
    defparam count_2226_add_4_10.INJECT1_0 = "NO";
    defparam count_2226_add_4_10.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_8 (.A0(\fcw_r[6] ), .B0(n184[6]), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[7] ), .B1(n184[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15764), .COUT(n15765), .S0(n124), .S1(n123));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_8.INIT0 = 16'h5666;
    defparam count_2226_add_4_8.INIT1 = 16'h5666;
    defparam count_2226_add_4_8.INJECT1_0 = "NO";
    defparam count_2226_add_4_8.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_6 (.A0(\fcw_r[4] ), .B0(n184[4]), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[5] ), .B1(n184[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15763), .COUT(n15764), .S0(n126), .S1(n125));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_6.INIT0 = 16'h5666;
    defparam count_2226_add_4_6.INIT1 = 16'h5666;
    defparam count_2226_add_4_6.INJECT1_0 = "NO";
    defparam count_2226_add_4_6.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_4 (.A0(\fcw_r[2] ), .B0(n184[2]), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[3] ), .B1(n184[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15762), .COUT(n15763), .S0(n128), .S1(n127));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_4.INIT0 = 16'h5666;
    defparam count_2226_add_4_4.INIT1 = 16'h5666;
    defparam count_2226_add_4_4.INJECT1_0 = "NO";
    defparam count_2226_add_4_4.INJECT1_1 = "NO";
    CCU2D count_2226_add_4_2 (.A0(\fcw_r[0] ), .B0(n25), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[1] ), .B1(n184[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15762), .S1(n129));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226_add_4_2.INIT0 = 16'h7000;
    defparam count_2226_add_4_2.INIT1 = 16'h5666;
    defparam count_2226_add_4_2.INJECT1_0 = "NO";
    defparam count_2226_add_4_2.INJECT1_1 = "NO";
    CCU2D add_4165_10 (.A0(yinjie[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15512), 
          .S1(n7621));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_4165_10.INIT0 = 16'h5aaa;
    defparam add_4165_10.INIT1 = 16'h0000;
    defparam add_4165_10.INJECT1_0 = "NO";
    defparam add_4165_10.INJECT1_1 = "NO";
    CCU2D add_4165_8 (.A0(yinjie[0]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(yinjie[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15511), .COUT(n15512));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_4165_8.INIT0 = 16'h5aaa;
    defparam add_4165_8.INIT1 = 16'h5aaa;
    defparam add_4165_8.INJECT1_0 = "NO";
    defparam add_4165_8.INJECT1_1 = "NO";
    CCU2D add_4165_6 (.A0(yinjie[2]), .B0(n8), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15510), 
          .COUT(n15511), .S0(n7610[5]), .S1(n7610[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_4165_6.INIT0 = 16'h7888;
    defparam add_4165_6.INIT1 = 16'hf000;
    defparam add_4165_6.INJECT1_0 = "NO";
    defparam add_4165_6.INJECT1_1 = "NO";
    CCU2D add_4165_4 (.A0(yinjie[2]), .B0(n9471), .C0(GND_net), .D0(GND_net), 
          .A1(yinjie[2]), .B1(n8), .C1(GND_net), .D1(GND_net), .CIN(n15509), 
          .COUT(n15510), .S0(n7610[3]), .S1(n7610[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_4165_4.INIT0 = 16'h9666;
    defparam add_4165_4.INIT1 = 16'h9666;
    defparam add_4165_4.INJECT1_0 = "NO";
    defparam add_4165_4.INJECT1_1 = "NO";
    CCU2D add_4165_2 (.A0(yinjie[1]), .B0(yinjie[0]), .C0(GND_net), .D0(GND_net), 
          .A1(yinjie[1]), .B1(yinjie[0]), .C1(yinjie[2]), .D1(GND_net), 
          .COUT(n15509), .S1(n7610[2]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_4165_2.INIT0 = 16'h7000;
    defparam add_4165_2.INIT1 = 16'h9696;
    defparam add_4165_2.INJECT1_0 = "NO";
    defparam add_4165_2.INJECT1_1 = "NO";
    LUT4 i15_4_lut (.A(n7597[5]), .B(\yinjie_box[1] ), .C(n19846), .D(\fcw_r_15__N_527[0] ), 
         .Z(fcw_r_15__N_527[5])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i15_4_lut.init = 16'hfaca;
    FD1S3DX count_2226__i0 (.D(n132[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n25)) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i0.GSR = "DISABLED";
    LUT4 i10511_4_lut_4_lut_4_lut (.A(\yinjie_box[1] ), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .D(n7597[8]), .Z(fcw_r_15__N_527[8])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i10511_4_lut_4_lut_4_lut.init = 16'h2f20;
    LUT4 i10474_3_lut_then_4_lut (.A(\fcw_r_15__N_527[0] ), .B(n19846), 
         .C(n7610[4]), .D(\yinjie_box[1] ), .Z(n18861)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (B+(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i10474_3_lut_then_4_lut.init = 16'h038b;
    LUT4 i10474_3_lut_else_4_lut (.A(\fcw_r_15__N_527[0] ), .B(n19846), 
         .C(n7610[4]), .D(\yinjie_box[1] ), .Z(n18860)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B+!(C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i10474_3_lut_else_4_lut.init = 16'h30b8;
    FD1S3AX fcw_r_i2 (.D(fcw_r_15__N_495[1]), .CK(clk_N_168), .Q(\fcw_r[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(fcw_r_15__N_495[2]), .CK(clk_N_168), .Q(\fcw_r[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_i4 (.D(fcw_r_15__N_495[3]), .CK(clk_N_168), .Q(\fcw_r[3] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_i5 (.D(fcw_r_15__N_527[4]), .CK(clk_N_168), .Q(\fcw_r[4] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_i6 (.D(fcw_r_15__N_527[5]), .CK(clk_N_168), .Q(\fcw_r[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_i7 (.D(fcw_r_15__N_527[6]), .CK(clk_N_168), .Q(\fcw_r[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_i8 (.D(fcw_r_15__N_527[7]), .CK(clk_N_168), .Q(\fcw_r[7] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i8.GSR = "DISABLED";
    FD1S3AX fcw_r_i9 (.D(fcw_r_15__N_527[8]), .CK(clk_N_168), .Q(\fcw_r[8] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i9.GSR = "DISABLED";
    FD1S3AX fcw_r_i10 (.D(fcw_r_15__N_495[9]), .CK(clk_N_168), .Q(\fcw_r[9] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i10.GSR = "DISABLED";
    FD1S3IX fcw_r_i11 (.D(n7597[10]), .CK(clk_N_168), .CD(stat), .Q(\fcw_r[10] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=47, LSE_RLINE=56 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i11.GSR = "DISABLED";
    LUT4 mux_1493_i1_3_lut_rep_603 (.A(yinjie[0]), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .Z(n18785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam mux_1493_i1_3_lut_rep_603.init = 16'hcaca;
    LUT4 i3589_2_lut_3_lut_4_lut (.A(yinjie[0]), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .D(yinjie[2]), .Z(\fcw_r_15__N_495[8] )) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3589_2_lut_3_lut_4_lut.init = 16'hc5ca;
    FD1S3DX count_2226__i1 (.D(n132[1]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i1.GSR = "DISABLED";
    FD1S3DX count_2226__i2 (.D(n132[2]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i2.GSR = "DISABLED";
    FD1S3DX count_2226__i3 (.D(n132[3]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i3.GSR = "DISABLED";
    FD1S3DX count_2226__i4 (.D(n132[4]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i4.GSR = "DISABLED";
    FD1S3DX count_2226__i5 (.D(n132[5]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i5.GSR = "DISABLED";
    FD1S3DX count_2226__i6 (.D(n132[6]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i6.GSR = "DISABLED";
    FD1S3DX count_2226__i7 (.D(n132[7]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i7.GSR = "DISABLED";
    FD1S3DX count_2226__i8 (.D(n132[8]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i8.GSR = "DISABLED";
    FD1S3DX count_2226__i9 (.D(n132[9]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i9.GSR = "DISABLED";
    FD1S3DX count_2226__i10 (.D(n132[10]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i10.GSR = "DISABLED";
    FD1S3DX count_2226__i11 (.D(n132[11]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i11.GSR = "DISABLED";
    FD1S3DX count_2226__i12 (.D(n132[12]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i12.GSR = "DISABLED";
    FD1S3DX count_2226__i13 (.D(n132[13]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(n184[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i13.GSR = "DISABLED";
    FD1S3DX count_2226__i14 (.D(n132[14]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[14] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i14.GSR = "DISABLED";
    FD1S3DX count_2226__i15 (.D(n132[15]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[15] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i15.GSR = "DISABLED";
    FD1S3DX count_2226__i16 (.D(n132[16]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[16] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i16.GSR = "DISABLED";
    FD1S3DX count_2226__i17 (.D(n132[17]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[17] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i17.GSR = "DISABLED";
    FD1S3DX count_2226__i18 (.D(n132[18]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[18] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i18.GSR = "DISABLED";
    FD1S3DX count_2226__i19 (.D(n132[19]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[19] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i19.GSR = "DISABLED";
    FD1S3DX count_2226__i20 (.D(n132[20]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[20] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i20.GSR = "DISABLED";
    FD1S3DX count_2226__i21 (.D(n132[21]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[21] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i21.GSR = "DISABLED";
    FD1S3DX count_2226__i22 (.D(n132[22]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[22] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i22.GSR = "DISABLED";
    FD1S3DX count_2226__i23 (.D(n132[23]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[23] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i23.GSR = "DISABLED";
    FD1S3DX count_2226__i24 (.D(n132[24]), .CK(clk__inv), .CD(pwm_out2_N_125), 
            .Q(\count1[24] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2226__i24.GSR = "DISABLED";
    CCU2D add_2977_8 (.A0(n7621), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15802), 
          .S0(n7597[10]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_2977_8.INIT0 = 16'h5aaa;
    defparam add_2977_8.INIT1 = 16'h0000;
    defparam add_2977_8.INJECT1_0 = "NO";
    defparam add_2977_8.INJECT1_1 = "NO";
    CCU2D add_2977_6 (.A0(yinjie[2]), .B0(n8), .C0(yinjie[1]), .D0(GND_net), 
          .A1(yinjie[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15801), .COUT(n15802), .S0(n7597[8]), .S1(n7597[9]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_2977_6.INIT0 = 16'h7878;
    defparam add_2977_6.INIT1 = 16'h5aaa;
    defparam add_2977_6.INJECT1_0 = "NO";
    defparam add_2977_6.INJECT1_1 = "NO";
    CCU2D add_2977_4 (.A0(n7610[6]), .B0(yinjie[1]), .C0(yinjie[2]), .D0(yinjie[0]), 
          .A1(yinjie[2]), .B1(n8), .C1(yinjie[0]), .D1(GND_net), .CIN(n15800), 
          .COUT(n15801), .S0(n7597[6]), .S1(n7597[7]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_2977_4.INIT0 = 16'h5a96;
    defparam add_2977_4.INIT1 = 16'h9696;
    defparam add_2977_4.INJECT1_0 = "NO";
    defparam add_2977_4.INJECT1_1 = "NO";
    LUT4 i2_2_lut_4_lut_4_lut_4_lut (.A(\yinjie_box[1] ), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .D(n7597[7]), .Z(fcw_r_15__N_527[7])) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i2_2_lut_4_lut_4_lut_4_lut.init = 16'h4f40;
    LUT4 mux_1493_i3_4_lut_4_lut (.A(\yinjie_box[1] ), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .D(n7610[2]), .Z(fcw_r_15__N_495[2])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam mux_1493_i3_4_lut_4_lut.init = 16'hefe0;
    LUT4 mux_1493_i4_3_lut_4_lut (.A(\yinjie_box[1] ), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .D(n7610[3]), .Z(fcw_r_15__N_495[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam mux_1493_i4_3_lut_4_lut.init = 16'h2f20;
    LUT4 i12_3_lut_4_lut (.A(\yinjie_box[1] ), .B(\fcw_r_15__N_527[0] ), 
         .C(n19846), .D(n7597[6]), .Z(fcw_r_15__N_527[6])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i12_3_lut_4_lut.init = 16'h2f20;
    CCU2D add_2977_2 (.A0(n7610[4]), .B0(yinjie[0]), .C0(GND_net), .D0(GND_net), 
          .A1(yinjie[1]), .B1(yinjie[0]), .C1(n7610[5]), .D1(GND_net), 
          .COUT(n15800), .S1(n7597[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam add_2977_2.INIT0 = 16'h7000;
    defparam add_2977_2.INIT1 = 16'h9696;
    defparam add_2977_2.INJECT1_0 = "NO";
    defparam add_2977_2.INJECT1_1 = "NO";
    LUT4 i5221_3_lut (.A(yinjie[1]), .B(yinjie[2]), .C(yinjie[0]), .Z(n8)) /* synthesis lut_function=(A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam i5221_3_lut.init = 16'ha8a8;
    LUT4 i4669_2_lut (.A(yinjie[1]), .B(yinjie[0]), .Z(n9471)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(17[17:27])
    defparam i4669_2_lut.init = 16'h2222;
    PFUMX i12630 (.BLUT(n18860), .ALUT(n18861), .C0(yinjie[0]), .Z(fcw_r_15__N_527[4]));
    LUT4 n7599_bdd_4_lut (.A(n7597[9]), .B(\yinjie_box[1] ), .C(n19846), 
         .D(\fcw_r_15__N_527[0] ), .Z(fcw_r_15__N_495[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam n7599_bdd_4_lut.init = 16'hca0a;
    LUT4 i10386_2_lut (.A(\yinjie_box[1] ), .B(\fcw_r_15__N_527[0] ), .Z(fcw_r_15__N_527[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(19[17:31])
    defparam i10386_2_lut.init = 16'h6666;
    LUT4 i10528_2_lut (.A(yinjie[1]), .B(yinjie[0]), .Z(n7610[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i10528_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module DDS_U8
//

module DDS_U8 (\count13[23] , GND_net, \count13[24] , \count_24__N_543[23] , 
            \count_24__N_543[24] , \count13[21] , \count13[22] , \count_24__N_543[21] , 
            \count_24__N_543[22] , \count13[19] , \count13[20] , \count_24__N_543[19] , 
            \count_24__N_543[20] , \count13[17] , \count13[18] , \count_24__N_543[17] , 
            \count_24__N_543[18] , \count13[15] , \count13[16] , \count_24__N_543[15] , 
            \count_24__N_543[16] , \count13[14] , \count_24__N_543[13] , 
            \count_24__N_543[14] , \fcw_r[10] , \count_24__N_543[11] , 
            \count_24__N_543[12] , \fcw_r[8] , \fcw_r[9] , \count_24__N_543[9] , 
            \count_24__N_543[10] , \fcw_r[6] , \fcw_r[7] , \count_24__N_543[7] , 
            \count_24__N_543[8] , \fcw_r[4] , \fcw_r[5] , \count_24__N_543[5] , 
            \count_24__N_543[6] , \fcw_r[2] , \fcw_r[3] , \count_24__N_543[3] , 
            \count_24__N_543[4] , \count13[1] , \fcw_r[0] , \fcw_r[1] , 
            \count_24__N_543[2] , clk, clk__inv, rst_n_c, key_pa_c, 
            pwm_out2_N_125, clk_N_168, n49, n48, n47, n46, n45, 
            n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
            n34, n33, n32, n31, n30, n29, n28, n27, n26) /* synthesis syn_module_defined=1 */ ;
    output \count13[23] ;
    input GND_net;
    output \count13[24] ;
    output \count_24__N_543[23] ;
    output \count_24__N_543[24] ;
    output \count13[21] ;
    output \count13[22] ;
    output \count_24__N_543[21] ;
    output \count_24__N_543[22] ;
    output \count13[19] ;
    output \count13[20] ;
    output \count_24__N_543[19] ;
    output \count_24__N_543[20] ;
    output \count13[17] ;
    output \count13[18] ;
    output \count_24__N_543[17] ;
    output \count_24__N_543[18] ;
    output \count13[15] ;
    output \count13[16] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[16] ;
    output \count13[14] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[14] ;
    input \fcw_r[10] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[12] ;
    input \fcw_r[8] ;
    input \fcw_r[9] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[10] ;
    input \fcw_r[6] ;
    input \fcw_r[7] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[8] ;
    input \fcw_r[4] ;
    input \fcw_r[5] ;
    output \count_24__N_543[5] ;
    output \count_24__N_543[6] ;
    input \fcw_r[2] ;
    input \fcw_r[3] ;
    output \count_24__N_543[3] ;
    output \count_24__N_543[4] ;
    output \count13[1] ;
    input \fcw_r[0] ;
    input \fcw_r[1] ;
    output \count_24__N_543[2] ;
    input clk;
    output clk__inv;
    input rst_n_c;
    input key_pa_c;
    output pwm_out2_N_125;
    input clk_N_168;
    input n49;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    
    wire clk /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15474, n15473, n15472, n15471, n15470, n15469;
    wire [24:0]count13;   // d:/fpga_project/lattice_diamond/piano/speaker.v(15[14:21])
    
    wire n15468, n15467, n15466, n15465, n15464;
    
    CCU2D add_2218_24 (.A0(\count13[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count13[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15474), .S0(\count_24__N_543[23] ), .S1(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_24.INIT0 = 16'h5aaa;
    defparam add_2218_24.INIT1 = 16'h5aaa;
    defparam add_2218_24.INJECT1_0 = "NO";
    defparam add_2218_24.INJECT1_1 = "NO";
    CCU2D add_2218_22 (.A0(\count13[21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count13[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15473), .COUT(n15474), .S0(\count_24__N_543[21] ), 
          .S1(\count_24__N_543[22] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_22.INIT0 = 16'h5aaa;
    defparam add_2218_22.INIT1 = 16'h5aaa;
    defparam add_2218_22.INJECT1_0 = "NO";
    defparam add_2218_22.INJECT1_1 = "NO";
    CCU2D add_2218_20 (.A0(\count13[19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count13[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15472), .COUT(n15473), .S0(\count_24__N_543[19] ), 
          .S1(\count_24__N_543[20] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_20.INIT0 = 16'h5aaa;
    defparam add_2218_20.INIT1 = 16'h5aaa;
    defparam add_2218_20.INJECT1_0 = "NO";
    defparam add_2218_20.INJECT1_1 = "NO";
    CCU2D add_2218_18 (.A0(\count13[17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count13[18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15471), .COUT(n15472), .S0(\count_24__N_543[17] ), 
          .S1(\count_24__N_543[18] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_18.INIT0 = 16'h5aaa;
    defparam add_2218_18.INIT1 = 16'h5aaa;
    defparam add_2218_18.INJECT1_0 = "NO";
    defparam add_2218_18.INJECT1_1 = "NO";
    CCU2D add_2218_16 (.A0(\count13[15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count13[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15470), .COUT(n15471), .S0(\count_24__N_543[15] ), 
          .S1(\count_24__N_543[16] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_16.INIT0 = 16'h5aaa;
    defparam add_2218_16.INIT1 = 16'h5aaa;
    defparam add_2218_16.INJECT1_0 = "NO";
    defparam add_2218_16.INJECT1_1 = "NO";
    CCU2D add_2218_14 (.A0(count13[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count13[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15469), .COUT(n15470), .S0(\count_24__N_543[13] ), .S1(\count_24__N_543[14] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_14.INIT0 = 16'h5aaa;
    defparam add_2218_14.INIT1 = 16'h5aaa;
    defparam add_2218_14.INJECT1_0 = "NO";
    defparam add_2218_14.INJECT1_1 = "NO";
    CCU2D add_2218_12 (.A0(count13[11]), .B0(\fcw_r[10] ), .C0(GND_net), 
          .D0(GND_net), .A1(count13[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15468), .COUT(n15469), .S0(\count_24__N_543[11] ), 
          .S1(\count_24__N_543[12] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_12.INIT0 = 16'h5666;
    defparam add_2218_12.INIT1 = 16'h5aaa;
    defparam add_2218_12.INJECT1_0 = "NO";
    defparam add_2218_12.INJECT1_1 = "NO";
    CCU2D add_2218_10 (.A0(count13[9]), .B0(\fcw_r[8] ), .C0(GND_net), 
          .D0(GND_net), .A1(count13[10]), .B1(\fcw_r[9] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n15467), .COUT(n15468), .S0(\count_24__N_543[9] ), 
          .S1(\count_24__N_543[10] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_10.INIT0 = 16'h5666;
    defparam add_2218_10.INIT1 = 16'h5666;
    defparam add_2218_10.INJECT1_0 = "NO";
    defparam add_2218_10.INJECT1_1 = "NO";
    CCU2D add_2218_8 (.A0(count13[7]), .B0(\fcw_r[6] ), .C0(GND_net), 
          .D0(GND_net), .A1(count13[8]), .B1(\fcw_r[7] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n15466), .COUT(n15467), .S0(\count_24__N_543[7] ), 
          .S1(\count_24__N_543[8] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_8.INIT0 = 16'h5666;
    defparam add_2218_8.INIT1 = 16'h5666;
    defparam add_2218_8.INJECT1_0 = "NO";
    defparam add_2218_8.INJECT1_1 = "NO";
    CCU2D add_2218_6 (.A0(count13[5]), .B0(\fcw_r[4] ), .C0(GND_net), 
          .D0(GND_net), .A1(count13[6]), .B1(\fcw_r[5] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n15465), .COUT(n15466), .S0(\count_24__N_543[5] ), 
          .S1(\count_24__N_543[6] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_6.INIT0 = 16'h5666;
    defparam add_2218_6.INIT1 = 16'h5666;
    defparam add_2218_6.INJECT1_0 = "NO";
    defparam add_2218_6.INJECT1_1 = "NO";
    CCU2D add_2218_4 (.A0(count13[3]), .B0(\fcw_r[2] ), .C0(GND_net), 
          .D0(GND_net), .A1(count13[4]), .B1(\fcw_r[3] ), .C1(GND_net), 
          .D1(GND_net), .CIN(n15464), .COUT(n15465), .S0(\count_24__N_543[3] ), 
          .S1(\count_24__N_543[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_4.INIT0 = 16'h5666;
    defparam add_2218_4.INIT1 = 16'h5666;
    defparam add_2218_4.INJECT1_0 = "NO";
    defparam add_2218_4.INJECT1_1 = "NO";
    CCU2D add_2218_2 (.A0(\count13[1] ), .B0(\fcw_r[0] ), .C0(GND_net), 
          .D0(GND_net), .A1(count13[2]), .B1(\fcw_r[1] ), .C1(GND_net), 
          .D1(GND_net), .COUT(n15464), .S1(\count_24__N_543[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2218_2.INIT0 = 16'h7000;
    defparam add_2218_2.INIT1 = 16'h5666;
    defparam add_2218_2.INJECT1_0 = "NO";
    defparam add_2218_2.INJECT1_1 = "NO";
    LUT4 clk_I_0_1_lut_rep_638 (.A(clk), .Z(clk__inv)) /* synthesis lut_function=(!(A)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(541[12:23])
    defparam clk_I_0_1_lut_rep_638.init = 16'h5555;
    LUT4 i12279_2_lut (.A(rst_n_c), .B(key_pa_c), .Z(pwm_out2_N_125)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(543[7:13])
    defparam i12279_2_lut.init = 16'h7777;
    FD1S3DX count__i1 (.D(n49), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count13[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i1.GSR = "DISABLED";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count13[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count13[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count13[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count13[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count13[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count13[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=188 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U9
//

module DDS_U9 (\count12[24] , GND_net, n106, \count12[22] , \count12[23] , 
            n108, n107, \count12[20] , \count12[21] , n110, n109, 
            \count12[18] , \count12[19] , n112, n111, \count12[16] , 
            \count12[17] , n114, n113, \count12[14] , \count12[15] , 
            n116, n115, n118, n117, \fcw_r[2] , n120, n119, \fcw_r[0] , 
            \fcw_r[1] , n122, n121, n124, n123, n126, n125, n128, 
            n127, n25, n129, clk_N_168, pwm_out2_N_125, n132, n18757, 
            \fcw_r_15__N_495[11] , yinjie, n18785, n18784, n19846, 
            \yinjie_box[1] , \fcw_r_15__N_527[0] ) /* synthesis syn_module_defined=1 */ ;
    output \count12[24] ;
    input GND_net;
    output n106;
    output \count12[22] ;
    output \count12[23] ;
    output n108;
    output n107;
    output \count12[20] ;
    output \count12[21] ;
    output n110;
    output n109;
    output \count12[18] ;
    output \count12[19] ;
    output n112;
    output n111;
    output \count12[16] ;
    output \count12[17] ;
    output n114;
    output n113;
    output \count12[14] ;
    output \count12[15] ;
    output n116;
    output n115;
    output n118;
    output n117;
    input \fcw_r[2] ;
    output n120;
    output n119;
    input \fcw_r[0] ;
    input \fcw_r[1] ;
    output n122;
    output n121;
    output n124;
    output n123;
    output n126;
    output n125;
    output n128;
    output n127;
    output n25;
    output n129;
    input clk_N_168;
    input pwm_out2_N_125;
    input [24:0]n132;
    input n18757;
    input \fcw_r_15__N_495[11] ;
    input [2:0]yinjie;
    input n18785;
    input n18784;
    input n19846;
    input \yinjie_box[1] ;
    input \fcw_r_15__N_527[0] ;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15721, n15720, n15719, n15718, n15717, n15716, n15715;
    wire [24:0]n184;
    
    wire n15714, n4, n18701;
    wire [12:0]n6813;
    
    wire n15713, n4_adj_832, n15712;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15711, n15710, n18776, n15805;
    wire [9:0]n8492;
    
    wire n8503, n15804, n15803;
    
    CCU2D count_2230_add_4_26 (.A0(\count12[24] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15721), .S0(n106));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_26.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_26.INIT1 = 16'h0000;
    defparam count_2230_add_4_26.INJECT1_0 = "NO";
    defparam count_2230_add_4_26.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_24 (.A0(\count12[22] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count12[23] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15720), .COUT(n15721), .S0(n108), .S1(n107));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_24.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_24.INIT1 = 16'hfaaa;
    defparam count_2230_add_4_24.INJECT1_0 = "NO";
    defparam count_2230_add_4_24.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_22 (.A0(\count12[20] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count12[21] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15719), .COUT(n15720), .S0(n110), .S1(n109));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_22.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_22.INIT1 = 16'hfaaa;
    defparam count_2230_add_4_22.INJECT1_0 = "NO";
    defparam count_2230_add_4_22.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_20 (.A0(\count12[18] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count12[19] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15718), .COUT(n15719), .S0(n112), .S1(n111));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_20.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_20.INIT1 = 16'hfaaa;
    defparam count_2230_add_4_20.INJECT1_0 = "NO";
    defparam count_2230_add_4_20.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_18 (.A0(\count12[16] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count12[17] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15717), .COUT(n15718), .S0(n114), .S1(n113));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_18.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_18.INIT1 = 16'hfaaa;
    defparam count_2230_add_4_18.INJECT1_0 = "NO";
    defparam count_2230_add_4_18.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_16 (.A0(\count12[14] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count12[15] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15716), .COUT(n15717), .S0(n116), .S1(n115));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_16.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_16.INIT1 = 16'hfaaa;
    defparam count_2230_add_4_16.INJECT1_0 = "NO";
    defparam count_2230_add_4_16.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_14 (.A0(n184[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n184[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15715), .COUT(n15716), .S0(n118), .S1(n117));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_14.INIT0 = 16'hfaaa;
    defparam count_2230_add_4_14.INIT1 = 16'hfaaa;
    defparam count_2230_add_4_14.INJECT1_0 = "NO";
    defparam count_2230_add_4_14.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_12 (.A0(\fcw_r[2] ), .B0(n4), .C0(n184[10]), 
          .D0(GND_net), .A1(n184[11]), .B1(n18701), .C1(\fcw_r[2] ), 
          .D1(n6813[10]), .CIN(n15714), .COUT(n15715), .S0(n120), .S1(n119));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_12.INIT0 = 16'h9696;
    defparam count_2230_add_4_12.INIT1 = 16'h566a;
    defparam count_2230_add_4_12.INJECT1_0 = "NO";
    defparam count_2230_add_4_12.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_10 (.A0(n6813[8]), .B0(\fcw_r[0] ), .C0(n184[8]), 
          .D0(GND_net), .A1(\fcw_r[1] ), .B1(n4_adj_832), .C1(n184[9]), 
          .D1(GND_net), .CIN(n15713), .COUT(n15714), .S0(n122), .S1(n121));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_10.INIT0 = 16'h9696;
    defparam count_2230_add_4_10.INIT1 = 16'h9696;
    defparam count_2230_add_4_10.INJECT1_0 = "NO";
    defparam count_2230_add_4_10.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_8 (.A0(fcw_r[6]), .B0(n184[6]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[7]), .B1(n184[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15712), .COUT(n15713), .S0(n124), .S1(n123));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_8.INIT0 = 16'h5666;
    defparam count_2230_add_4_8.INIT1 = 16'h5666;
    defparam count_2230_add_4_8.INJECT1_0 = "NO";
    defparam count_2230_add_4_8.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_6 (.A0(fcw_r[4]), .B0(n184[4]), .C0(GND_net), 
          .D0(GND_net), .A1(fcw_r[5]), .B1(n184[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15711), .COUT(n15712), .S0(n126), .S1(n125));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_6.INIT0 = 16'h5666;
    defparam count_2230_add_4_6.INIT1 = 16'h5666;
    defparam count_2230_add_4_6.INJECT1_0 = "NO";
    defparam count_2230_add_4_6.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_4 (.A0(\fcw_r[2] ), .B0(n184[2]), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[0] ), .B1(n184[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n15710), .COUT(n15711), .S0(n128), .S1(n127));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_4.INIT0 = 16'h5666;
    defparam count_2230_add_4_4.INIT1 = 16'h5666;
    defparam count_2230_add_4_4.INJECT1_0 = "NO";
    defparam count_2230_add_4_4.INJECT1_1 = "NO";
    CCU2D count_2230_add_4_2 (.A0(\fcw_r[0] ), .B0(n25), .C0(GND_net), 
          .D0(GND_net), .A1(\fcw_r[1] ), .B1(n184[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15710), .S1(n129));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230_add_4_2.INIT0 = 16'h7000;
    defparam count_2230_add_4_2.INIT1 = 16'h5666;
    defparam count_2230_add_4_2.INJECT1_0 = "NO";
    defparam count_2230_add_4_2.INJECT1_1 = "NO";
    FD1S3DX count_2230__i0 (.D(n132[0]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n25)) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(\fcw_r[1] ), .B(n18776), .C(n6813[9]), .D(n6813[10]), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_4_lut.init = 16'h17e8;
    LUT4 i3846_2_lut_rep_594 (.A(n6813[8]), .B(\fcw_r[0] ), .Z(n18776)) /* synthesis lut_function=(A (B)) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3846_2_lut_rep_594.init = 16'h8888;
    LUT4 i3857_4_lut_3_lut_rep_519_4_lut (.A(n6813[8]), .B(\fcw_r[0] ), 
         .C(n6813[9]), .D(\fcw_r[1] ), .Z(n18701)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i3857_4_lut_3_lut_rep_519_4_lut.init = 16'hf880;
    LUT4 i1_2_lut_3_lut (.A(n6813[8]), .B(\fcw_r[0] ), .C(n6813[9]), .Z(n4_adj_832)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    CCU2D add_3786_7 (.A0(n18757), .B0(\fcw_r_15__N_495[11] ), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15805), .S0(n8492[9]), .S1(n8503));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3786_7.INIT0 = 16'h7888;
    defparam add_3786_7.INIT1 = 16'h0000;
    defparam add_3786_7.INJECT1_0 = "NO";
    defparam add_3786_7.INJECT1_1 = "NO";
    FD1S3AX fcw_r_ret0_i4 (.D(n8492[4]), .CK(clk_N_168), .Q(fcw_r[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_ret0_i5 (.D(n8492[5]), .CK(clk_N_168), .Q(fcw_r[5]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_ret0_i6 (.D(n8492[6]), .CK(clk_N_168), .Q(fcw_r[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_ret0_i7 (.D(n8492[7]), .CK(clk_N_168), .Q(fcw_r[7]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_ret0_i8 (.D(n8492[8]), .CK(clk_N_168), .Q(n6813[8]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i8.GSR = "DISABLED";
    FD1S3AX fcw_r_ret0_i9 (.D(n8492[9]), .CK(clk_N_168), .Q(n6813[9]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i9.GSR = "DISABLED";
    FD1S3AX fcw_r_ret0_i10 (.D(n8503), .CK(clk_N_168), .Q(n6813[10]));   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_ret0_i10.GSR = "DISABLED";
    CCU2D add_3786_5 (.A0(yinjie[2]), .B0(n18785), .C0(n18784), .D0(n19846), 
          .A1(n18757), .B1(\fcw_r_15__N_495[11] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15804), .COUT(n15805), .S0(n8492[7]), .S1(n8492[8]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3786_5.INIT0 = 16'hf078;
    defparam add_3786_5.INIT1 = 16'h9666;
    defparam add_3786_5.INJECT1_0 = "NO";
    defparam add_3786_5.INJECT1_1 = "NO";
    CCU2D add_3786_3 (.A0(yinjie[2]), .B0(n19846), .C0(\yinjie_box[1] ), 
          .D0(yinjie[1]), .A1(yinjie[2]), .B1(yinjie[0]), .C1(\fcw_r_15__N_527[0] ), 
          .D1(n19846), .CIN(n15803), .COUT(n15804), .S0(n8492[5]), .S1(n8492[6]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3786_3.INIT0 = 16'hd1e2;
    defparam add_3786_3.INIT1 = 16'hf066;
    defparam add_3786_3.INJECT1_0 = "NO";
    defparam add_3786_3.INJECT1_1 = "NO";
    CCU2D add_3786_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n18784), .B1(n19846), .C1(\fcw_r_15__N_527[0] ), .D1(yinjie[0]), 
          .COUT(n15803), .S1(n8492[4]));   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam add_3786_1.INIT0 = 16'hF000;
    defparam add_3786_1.INIT1 = 16'h596a;
    defparam add_3786_1.INJECT1_0 = "NO";
    defparam add_3786_1.INJECT1_1 = "NO";
    FD1S3DX count_2230__i1 (.D(n132[1]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i1.GSR = "DISABLED";
    FD1S3DX count_2230__i2 (.D(n132[2]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i2.GSR = "DISABLED";
    FD1S3DX count_2230__i3 (.D(n132[3]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i3.GSR = "DISABLED";
    FD1S3DX count_2230__i4 (.D(n132[4]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i4.GSR = "DISABLED";
    FD1S3DX count_2230__i5 (.D(n132[5]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i5.GSR = "DISABLED";
    FD1S3DX count_2230__i6 (.D(n132[6]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i6.GSR = "DISABLED";
    FD1S3DX count_2230__i7 (.D(n132[7]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i7.GSR = "DISABLED";
    FD1S3DX count_2230__i8 (.D(n132[8]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i8.GSR = "DISABLED";
    FD1S3DX count_2230__i9 (.D(n132[9]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i9.GSR = "DISABLED";
    FD1S3DX count_2230__i10 (.D(n132[10]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i10.GSR = "DISABLED";
    FD1S3DX count_2230__i11 (.D(n132[11]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i11.GSR = "DISABLED";
    FD1S3DX count_2230__i12 (.D(n132[12]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i12.GSR = "DISABLED";
    FD1S3DX count_2230__i13 (.D(n132[13]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(n184[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i13.GSR = "DISABLED";
    FD1S3DX count_2230__i14 (.D(n132[14]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[14] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i14.GSR = "DISABLED";
    FD1S3DX count_2230__i15 (.D(n132[15]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[15] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i15.GSR = "DISABLED";
    FD1S3DX count_2230__i16 (.D(n132[16]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[16] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i16.GSR = "DISABLED";
    FD1S3DX count_2230__i17 (.D(n132[17]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[17] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i17.GSR = "DISABLED";
    FD1S3DX count_2230__i18 (.D(n132[18]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[18] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i18.GSR = "DISABLED";
    FD1S3DX count_2230__i19 (.D(n132[19]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[19] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i19.GSR = "DISABLED";
    FD1S3DX count_2230__i20 (.D(n132[20]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[20] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i20.GSR = "DISABLED";
    FD1S3DX count_2230__i21 (.D(n132[21]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[21] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i21.GSR = "DISABLED";
    FD1S3DX count_2230__i22 (.D(n132[22]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[22] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i22.GSR = "DISABLED";
    FD1S3DX count_2230__i23 (.D(n132[23]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[23] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i23.GSR = "DISABLED";
    FD1S3DX count_2230__i24 (.D(n132[24]), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count12[24] )) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam count_2230__i24.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U10
//

module DDS_U10 (clk_N_168, n18705, \count11[23] , GND_net, \count11[24] , 
            \count_24__N_543[23] , \count_24__N_543[24] , \count11[21] , 
            \count11[22] , \count_24__N_543[21] , \count_24__N_543[22] , 
            \count11[19] , \count11[20] , \count_24__N_543[19] , \count_24__N_543[20] , 
            \count11[17] , \count11[18] , \count_24__N_543[17] , \count_24__N_543[18] , 
            \count11[15] , \count11[16] , \count_24__N_543[15] , \count_24__N_543[16] , 
            \count11[14] , \count_24__N_543[13] , \count_24__N_543[14] , 
            \count_24__N_543[11] , \count_24__N_543[12] , \count_24__N_543[9] , 
            \count_24__N_543[10] , \count_24__N_543[7] , \count_24__N_543[8] , 
            \fcw_r[6] , \count_24__N_543[5] , \count_24__N_543[6] , \count_24__N_543[3] , 
            \count_24__N_543[4] , \count11[1] , \count_24__N_543[2] , 
            n18757, n18716, \fcw_r_15__N_495[11] , n18634, n18608, 
            pwm_out2_N_125, n49, n48, n47, n46, n45, n44, n43, 
            n42, n41, n40, n39, n38, n37, n36, n35, n34, n33, 
            n32, n31, n30, n29, n28, n27, n26, n18717, n19839, 
            n19840, n18785, n18784, \fcw_r_15__N_495[8] , \fcw_r_15__N_495[9] , 
            \fcw_r_15__N_495[10] ) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    input n18705;
    output \count11[23] ;
    input GND_net;
    output \count11[24] ;
    output \count_24__N_543[23] ;
    output \count_24__N_543[24] ;
    output \count11[21] ;
    output \count11[22] ;
    output \count_24__N_543[21] ;
    output \count_24__N_543[22] ;
    output \count11[19] ;
    output \count11[20] ;
    output \count_24__N_543[19] ;
    output \count_24__N_543[20] ;
    output \count11[17] ;
    output \count11[18] ;
    output \count_24__N_543[17] ;
    output \count_24__N_543[18] ;
    output \count11[15] ;
    output \count11[16] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[16] ;
    output \count11[14] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[14] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[12] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[10] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[8] ;
    output \fcw_r[6] ;
    output \count_24__N_543[5] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[3] ;
    output \count_24__N_543[4] ;
    output \count11[1] ;
    output \count_24__N_543[2] ;
    input n18757;
    input n18716;
    input \fcw_r_15__N_495[11] ;
    input n18634;
    output n18608;
    input pwm_out2_N_125;
    input n49;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    input n18717;
    input n19839;
    input n19840;
    input n18785;
    input n18784;
    input \fcw_r_15__N_495[8] ;
    input \fcw_r_15__N_495[9] ;
    input \fcw_r_15__N_495[10] ;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15454, n15453, n15452, n15451, n15450, n15449;
    wire [24:0]count11;   // d:/fpga_project/lattice_diamond/piano/speaker.v(14[34:41])
    
    wire n15448, n15447, n15446, n15445, n15444;
    
    FD1S3AX fcw_r_i1 (.D(n18705), .CK(clk_N_168), .Q(fcw_r[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D add_2214_24 (.A0(\count11[23] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count11[24] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15454), .S0(\count_24__N_543[23] ), .S1(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_24.INIT0 = 16'h5aaa;
    defparam add_2214_24.INIT1 = 16'h5aaa;
    defparam add_2214_24.INJECT1_0 = "NO";
    defparam add_2214_24.INJECT1_1 = "NO";
    CCU2D add_2214_22 (.A0(\count11[21] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count11[22] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15453), .COUT(n15454), .S0(\count_24__N_543[21] ), 
          .S1(\count_24__N_543[22] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_22.INIT0 = 16'h5aaa;
    defparam add_2214_22.INIT1 = 16'h5aaa;
    defparam add_2214_22.INJECT1_0 = "NO";
    defparam add_2214_22.INJECT1_1 = "NO";
    CCU2D add_2214_20 (.A0(\count11[19] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count11[20] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15452), .COUT(n15453), .S0(\count_24__N_543[19] ), 
          .S1(\count_24__N_543[20] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_20.INIT0 = 16'h5aaa;
    defparam add_2214_20.INIT1 = 16'h5aaa;
    defparam add_2214_20.INJECT1_0 = "NO";
    defparam add_2214_20.INJECT1_1 = "NO";
    CCU2D add_2214_18 (.A0(\count11[17] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count11[18] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15451), .COUT(n15452), .S0(\count_24__N_543[17] ), 
          .S1(\count_24__N_543[18] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_18.INIT0 = 16'h5aaa;
    defparam add_2214_18.INIT1 = 16'h5aaa;
    defparam add_2214_18.INJECT1_0 = "NO";
    defparam add_2214_18.INJECT1_1 = "NO";
    CCU2D add_2214_16 (.A0(\count11[15] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\count11[16] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15450), .COUT(n15451), .S0(\count_24__N_543[15] ), 
          .S1(\count_24__N_543[16] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_16.INIT0 = 16'h5aaa;
    defparam add_2214_16.INIT1 = 16'h5aaa;
    defparam add_2214_16.INJECT1_0 = "NO";
    defparam add_2214_16.INJECT1_1 = "NO";
    CCU2D add_2214_14 (.A0(count11[13]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count11[14] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15449), .COUT(n15450), .S0(\count_24__N_543[13] ), .S1(\count_24__N_543[14] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_14.INIT0 = 16'h5aaa;
    defparam add_2214_14.INIT1 = 16'h5aaa;
    defparam add_2214_14.INJECT1_0 = "NO";
    defparam add_2214_14.INJECT1_1 = "NO";
    CCU2D add_2214_12 (.A0(count11[11]), .B0(fcw_r[11]), .C0(GND_net), 
          .D0(GND_net), .A1(count11[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15448), .COUT(n15449), .S0(\count_24__N_543[11] ), 
          .S1(\count_24__N_543[12] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_12.INIT0 = 16'h5666;
    defparam add_2214_12.INIT1 = 16'h5aaa;
    defparam add_2214_12.INJECT1_0 = "NO";
    defparam add_2214_12.INJECT1_1 = "NO";
    CCU2D add_2214_10 (.A0(count11[9]), .B0(fcw_r[9]), .C0(GND_net), .D0(GND_net), 
          .A1(count11[10]), .B1(fcw_r[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15447), .COUT(n15448), .S0(\count_24__N_543[9] ), .S1(\count_24__N_543[10] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_10.INIT0 = 16'h5666;
    defparam add_2214_10.INIT1 = 16'h5666;
    defparam add_2214_10.INJECT1_0 = "NO";
    defparam add_2214_10.INJECT1_1 = "NO";
    CCU2D add_2214_8 (.A0(count11[7]), .B0(fcw_r[7]), .C0(GND_net), .D0(GND_net), 
          .A1(count11[8]), .B1(fcw_r[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15446), .COUT(n15447), .S0(\count_24__N_543[7] ), .S1(\count_24__N_543[8] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_8.INIT0 = 16'h5666;
    defparam add_2214_8.INIT1 = 16'h5666;
    defparam add_2214_8.INJECT1_0 = "NO";
    defparam add_2214_8.INJECT1_1 = "NO";
    CCU2D add_2214_6 (.A0(count11[5]), .B0(fcw_r[5]), .C0(GND_net), .D0(GND_net), 
          .A1(count11[6]), .B1(\fcw_r[6] ), .C1(GND_net), .D1(GND_net), 
          .CIN(n15445), .COUT(n15446), .S0(\count_24__N_543[5] ), .S1(\count_24__N_543[6] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_6.INIT0 = 16'h5666;
    defparam add_2214_6.INIT1 = 16'h5666;
    defparam add_2214_6.INJECT1_0 = "NO";
    defparam add_2214_6.INJECT1_1 = "NO";
    CCU2D add_2214_4 (.A0(count11[3]), .B0(fcw_r[3]), .C0(GND_net), .D0(GND_net), 
          .A1(count11[4]), .B1(fcw_r[4]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15444), .COUT(n15445), .S0(\count_24__N_543[3] ), .S1(\count_24__N_543[4] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_4.INIT0 = 16'h5666;
    defparam add_2214_4.INIT1 = 16'h5666;
    defparam add_2214_4.INJECT1_0 = "NO";
    defparam add_2214_4.INJECT1_1 = "NO";
    CCU2D add_2214_2 (.A0(\count11[1] ), .B0(\fcw_r[6] ), .C0(GND_net), 
          .D0(GND_net), .A1(count11[2]), .B1(fcw_r[2]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15444), .S1(\count_24__N_543[2] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_2214_2.INIT0 = 16'h7000;
    defparam add_2214_2.INIT1 = 16'h5666;
    defparam add_2214_2.INJECT1_0 = "NO";
    defparam add_2214_2.INJECT1_1 = "NO";
    LUT4 i4146_4_lut_3_lut_rep_426_4_lut (.A(n18757), .B(n18716), .C(\fcw_r_15__N_495[11] ), 
         .D(n18634), .Z(n18608)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i4146_4_lut_3_lut_rep_426_4_lut.init = 16'hf660;
    FD1S3DX count__i1 (.D(n49), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count11[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i1.GSR = "DISABLED";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count11[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count11[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count11[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count11[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count11[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count11[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    FD1S3AX fcw_r_i2 (.D(n18717), .CK(clk_N_168), .Q(fcw_r[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(n19839), .CK(clk_N_168), .Q(fcw_r[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_i4 (.D(n19840), .CK(clk_N_168), .Q(fcw_r[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_i5 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_i6 (.D(n18784), .CK(clk_N_168), .Q(fcw_r[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_i7 (.D(\fcw_r_15__N_495[8] ), .CK(clk_N_168), .Q(fcw_r[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_i8 (.D(\fcw_r_15__N_495[9] ), .CK(clk_N_168), .Q(fcw_r[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i8.GSR = "DISABLED";
    FD1S3AX fcw_r_i9 (.D(\fcw_r_15__N_495[10] ), .CK(clk_N_168), .Q(fcw_r[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i9.GSR = "DISABLED";
    FD1S3AX fcw_r_i10 (.D(\fcw_r_15__N_495[11] ), .CK(clk_N_168), .Q(fcw_r[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=157, LSE_RLINE=166 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i10.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module DDS_U11
//

module DDS_U11 (\fcw_r[2] , clk_N_168, n18785, \count10[24] , GND_net, 
            \count_24__N_543[24] , \count10[22] , \count10[23] , \count_24__N_543[22] , 
            \count_24__N_543[23] , \count10[20] , \count10[21] , \count_24__N_543[20] , 
            \count_24__N_543[21] , \count10[18] , \count10[19] , \count_24__N_543[18] , 
            \count_24__N_543[19] , \count10[16] , \count10[17] , \count_24__N_543[16] , 
            \count_24__N_543[17] , \count10[14] , \count10[15] , \count_24__N_543[14] , 
            \count_24__N_543[15] , \count_24__N_543[12] , \count_24__N_543[13] , 
            \count_24__N_543[10] , \count_24__N_543[11] , \count_24__N_543[8] , 
            \count_24__N_543[9] , \count_24__N_543[6] , \count_24__N_543[7] , 
            \count_24__N_543[4] , \count_24__N_543[5] , \count10[2] , 
            \count_24__N_543[3] , pwm_out2_N_125, n48, n47, n46, n45, 
            n44, n43, n42, n41, n40, n39, n38, n37, n36, n35, 
            n34, n33, n32, n31, n30, n29, n28, n27, n26, n18784, 
            \fcw_r_15__N_495[8] , \fcw_r_15__N_495[5] , \fcw_r_15__N_495[6] , 
            \fcw_r_15__N_495[8]_adj_10 , \fcw_r_15__N_495[9] , \fcw_r_15__N_495[10] , 
            n19846, \yinjie[2] , n18757, \fcw_r_15__N_495[11] , n18716, 
            n18634, n15966, n18690, n18705, n16936, n10972) /* synthesis syn_module_defined=1 */ ;
    output \fcw_r[2] ;
    input clk_N_168;
    input n18785;
    output \count10[24] ;
    input GND_net;
    output \count_24__N_543[24] ;
    output \count10[22] ;
    output \count10[23] ;
    output \count_24__N_543[22] ;
    output \count_24__N_543[23] ;
    output \count10[20] ;
    output \count10[21] ;
    output \count_24__N_543[20] ;
    output \count_24__N_543[21] ;
    output \count10[18] ;
    output \count10[19] ;
    output \count_24__N_543[18] ;
    output \count_24__N_543[19] ;
    output \count10[16] ;
    output \count10[17] ;
    output \count_24__N_543[16] ;
    output \count_24__N_543[17] ;
    output \count10[14] ;
    output \count10[15] ;
    output \count_24__N_543[14] ;
    output \count_24__N_543[15] ;
    output \count_24__N_543[12] ;
    output \count_24__N_543[13] ;
    output \count_24__N_543[10] ;
    output \count_24__N_543[11] ;
    output \count_24__N_543[8] ;
    output \count_24__N_543[9] ;
    output \count_24__N_543[6] ;
    output \count_24__N_543[7] ;
    output \count_24__N_543[4] ;
    output \count_24__N_543[5] ;
    output \count10[2] ;
    output \count_24__N_543[3] ;
    input pwm_out2_N_125;
    input n48;
    input n47;
    input n46;
    input n45;
    input n44;
    input n43;
    input n42;
    input n41;
    input n40;
    input n39;
    input n38;
    input n37;
    input n36;
    input n35;
    input n34;
    input n33;
    input n32;
    input n31;
    input n30;
    input n29;
    input n28;
    input n27;
    input n26;
    input n18784;
    input \fcw_r_15__N_495[8] ;
    input \fcw_r_15__N_495[5] ;
    input \fcw_r_15__N_495[6] ;
    input \fcw_r_15__N_495[8]_adj_10 ;
    input \fcw_r_15__N_495[9] ;
    input \fcw_r_15__N_495[10] ;
    input n19846;
    input \yinjie[2] ;
    input n18757;
    input \fcw_r_15__N_495[11] ;
    input n18716;
    output n18634;
    output n15966;
    input n18690;
    input n18705;
    output n16936;
    input n10972;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15442, n15441, n15440, n15439, n15438, n15437, n15436;
    wire [24:0]count10;   // d:/fpga_project/lattice_diamond/piano/speaker.v(14[14:21])
    
    wire n15435;
    wire [15:0]fcw_r;   // d:/fpga_project/lattice_diamond/piano/dds.v(12[13:18])
    
    wire n15434, n15433, n15432;
    wire [15:0]fcw_r_15__N_495;
    
    FD1S3AX fcw_r_i1 (.D(n18785), .CK(clk_N_168), .Q(\fcw_r[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i1.GSR = "DISABLED";
    CCU2D add_15_24 (.A0(\count10[24] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15442), 
          .S0(\count_24__N_543[24] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_24.INIT0 = 16'h5aaa;
    defparam add_15_24.INIT1 = 16'h0000;
    defparam add_15_24.INJECT1_0 = "NO";
    defparam add_15_24.INJECT1_1 = "NO";
    CCU2D add_15_22 (.A0(\count10[22] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count10[23] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15441), .COUT(n15442), .S0(\count_24__N_543[22] ), .S1(\count_24__N_543[23] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_22.INIT0 = 16'h5aaa;
    defparam add_15_22.INIT1 = 16'h5aaa;
    defparam add_15_22.INJECT1_0 = "NO";
    defparam add_15_22.INJECT1_1 = "NO";
    CCU2D add_15_20 (.A0(\count10[20] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count10[21] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15440), .COUT(n15441), .S0(\count_24__N_543[20] ), .S1(\count_24__N_543[21] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_20.INIT0 = 16'h5aaa;
    defparam add_15_20.INIT1 = 16'h5aaa;
    defparam add_15_20.INJECT1_0 = "NO";
    defparam add_15_20.INJECT1_1 = "NO";
    CCU2D add_15_18 (.A0(\count10[18] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count10[19] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15439), .COUT(n15440), .S0(\count_24__N_543[18] ), .S1(\count_24__N_543[19] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_18.INIT0 = 16'h5aaa;
    defparam add_15_18.INIT1 = 16'h5aaa;
    defparam add_15_18.INJECT1_0 = "NO";
    defparam add_15_18.INJECT1_1 = "NO";
    CCU2D add_15_16 (.A0(\count10[16] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count10[17] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15438), .COUT(n15439), .S0(\count_24__N_543[16] ), .S1(\count_24__N_543[17] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_16.INIT0 = 16'h5aaa;
    defparam add_15_16.INIT1 = 16'h5aaa;
    defparam add_15_16.INJECT1_0 = "NO";
    defparam add_15_16.INJECT1_1 = "NO";
    CCU2D add_15_14 (.A0(\count10[14] ), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\count10[15] ), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15437), .COUT(n15438), .S0(\count_24__N_543[14] ), .S1(\count_24__N_543[15] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_14.INIT0 = 16'h5aaa;
    defparam add_15_14.INIT1 = 16'h5aaa;
    defparam add_15_14.INJECT1_0 = "NO";
    defparam add_15_14.INJECT1_1 = "NO";
    CCU2D add_15_12 (.A0(count10[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count10[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15436), .COUT(n15437), .S0(\count_24__N_543[12] ), .S1(\count_24__N_543[13] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_12.INIT0 = 16'h5aaa;
    defparam add_15_12.INIT1 = 16'h5aaa;
    defparam add_15_12.INJECT1_0 = "NO";
    defparam add_15_12.INJECT1_1 = "NO";
    CCU2D add_15_10 (.A0(count10[10]), .B0(fcw_r[10]), .C0(GND_net), .D0(GND_net), 
          .A1(count10[11]), .B1(fcw_r[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15435), .COUT(n15436), .S0(\count_24__N_543[10] ), .S1(\count_24__N_543[11] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_10.INIT0 = 16'h5666;
    defparam add_15_10.INIT1 = 16'h5666;
    defparam add_15_10.INJECT1_0 = "NO";
    defparam add_15_10.INJECT1_1 = "NO";
    CCU2D add_15_8 (.A0(count10[8]), .B0(fcw_r[8]), .C0(GND_net), .D0(GND_net), 
          .A1(count10[9]), .B1(fcw_r[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15434), .COUT(n15435), .S0(\count_24__N_543[8] ), .S1(\count_24__N_543[9] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_8.INIT0 = 16'h5666;
    defparam add_15_8.INIT1 = 16'h5666;
    defparam add_15_8.INJECT1_0 = "NO";
    defparam add_15_8.INJECT1_1 = "NO";
    CCU2D add_15_6 (.A0(count10[6]), .B0(fcw_r[6]), .C0(GND_net), .D0(GND_net), 
          .A1(count10[7]), .B1(fcw_r[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15433), .COUT(n15434), .S0(\count_24__N_543[6] ), .S1(\count_24__N_543[7] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_6.INIT0 = 16'h5666;
    defparam add_15_6.INIT1 = 16'h5666;
    defparam add_15_6.INJECT1_0 = "NO";
    defparam add_15_6.INJECT1_1 = "NO";
    CCU2D add_15_4 (.A0(count10[4]), .B0(fcw_r[4]), .C0(GND_net), .D0(GND_net), 
          .A1(count10[5]), .B1(fcw_r[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n15432), .COUT(n15433), .S0(\count_24__N_543[4] ), .S1(\count_24__N_543[5] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_4.INIT0 = 16'h5666;
    defparam add_15_4.INIT1 = 16'h5666;
    defparam add_15_4.INJECT1_0 = "NO";
    defparam add_15_4.INJECT1_1 = "NO";
    CCU2D add_15_2 (.A0(\count10[2] ), .B0(\fcw_r[2] ), .C0(GND_net), 
          .D0(GND_net), .A1(count10[3]), .B1(fcw_r[3]), .C1(GND_net), 
          .D1(GND_net), .COUT(n15432), .S1(\count_24__N_543[3] ));   // d:/fpga_project/lattice_diamond/piano/dds.v(28[12:23])
    defparam add_15_2.INIT0 = 16'h7000;
    defparam add_15_2.INIT1 = 16'h5666;
    defparam add_15_2.INJECT1_0 = "NO";
    defparam add_15_2.INJECT1_1 = "NO";
    FD1S3DX count__i2 (.D(n48), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(\count10[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i2.GSR = "DISABLED";
    FD1S3DX count__i3 (.D(n47), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i3.GSR = "DISABLED";
    FD1S3DX count__i4 (.D(n46), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i4.GSR = "DISABLED";
    FD1S3DX count__i5 (.D(n45), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i5.GSR = "DISABLED";
    FD1S3DX count__i6 (.D(n44), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i6.GSR = "DISABLED";
    FD1S3DX count__i7 (.D(n43), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i7.GSR = "DISABLED";
    FD1S3DX count__i8 (.D(n42), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i8.GSR = "DISABLED";
    FD1S3DX count__i9 (.D(n41), .CK(clk_N_168), .CD(pwm_out2_N_125), .Q(count10[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i9.GSR = "DISABLED";
    FD1S3DX count__i10 (.D(n40), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count10[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i10.GSR = "DISABLED";
    FD1S3DX count__i11 (.D(n39), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count10[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i11.GSR = "DISABLED";
    FD1S3DX count__i12 (.D(n38), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count10[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i12.GSR = "DISABLED";
    FD1S3DX count__i13 (.D(n37), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(count10[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i13.GSR = "DISABLED";
    FD1S3DX count__i14 (.D(n36), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i14.GSR = "DISABLED";
    FD1S3DX count__i15 (.D(n35), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[15] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i15.GSR = "DISABLED";
    FD1S3DX count__i16 (.D(n34), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[16] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i16.GSR = "DISABLED";
    FD1S3DX count__i17 (.D(n33), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[17] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i17.GSR = "DISABLED";
    FD1S3DX count__i18 (.D(n32), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[18] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i18.GSR = "DISABLED";
    FD1S3DX count__i19 (.D(n31), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[19] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i19.GSR = "DISABLED";
    FD1S3DX count__i20 (.D(n30), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[20] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i20.GSR = "DISABLED";
    FD1S3DX count__i21 (.D(n29), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[21] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i21.GSR = "DISABLED";
    FD1S3DX count__i22 (.D(n28), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[22] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i22.GSR = "DISABLED";
    FD1S3DX count__i23 (.D(n27), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[23] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i23.GSR = "DISABLED";
    FD1S3DX count__i24 (.D(n26), .CK(clk_N_168), .CD(pwm_out2_N_125), 
            .Q(\count10[24] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(27[12] 30[16])
    defparam count__i24.GSR = "DISABLED";
    FD1S3AX fcw_r_i2 (.D(n18784), .CK(clk_N_168), .Q(fcw_r[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i2.GSR = "DISABLED";
    FD1S3AX fcw_r_i3 (.D(\fcw_r_15__N_495[8] ), .CK(clk_N_168), .Q(fcw_r[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i3.GSR = "DISABLED";
    FD1S3AX fcw_r_i4 (.D(\fcw_r_15__N_495[5] ), .CK(clk_N_168), .Q(fcw_r[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i4.GSR = "DISABLED";
    FD1S3AX fcw_r_i5 (.D(\fcw_r_15__N_495[6] ), .CK(clk_N_168), .Q(fcw_r[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i5.GSR = "DISABLED";
    FD1S3AX fcw_r_i6 (.D(fcw_r_15__N_495[7]), .CK(clk_N_168), .Q(fcw_r[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i6.GSR = "DISABLED";
    FD1S3AX fcw_r_i7 (.D(\fcw_r_15__N_495[8]_adj_10 ), .CK(clk_N_168), .Q(fcw_r[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i7.GSR = "DISABLED";
    FD1S3AX fcw_r_i8 (.D(\fcw_r_15__N_495[9] ), .CK(clk_N_168), .Q(fcw_r[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i8.GSR = "DISABLED";
    FD1S3AX fcw_r_i9 (.D(\fcw_r_15__N_495[10] ), .CK(clk_N_168), .Q(fcw_r[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i9.GSR = "DISABLED";
    LUT4 n18784_bdd_4_lut (.A(n18784), .B(n18785), .C(n19846), .D(\yinjie[2] ), 
         .Z(fcw_r_15__N_495[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam n18784_bdd_4_lut.init = 16'h8188;
    LUT4 i2_3_lut_4_lut (.A(n18757), .B(\fcw_r_15__N_495[11] ), .C(n18716), 
         .D(n18634), .Z(n15966)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i2_3_lut_4_lut.init = 16'h2dd2;
    LUT4 i4139_4_lut_3_lut_rep_452_4_lut (.A(n18757), .B(\fcw_r_15__N_495[11] ), 
         .C(n18690), .D(n18705), .Z(n18634)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i4139_4_lut_3_lut_rep_452_4_lut.init = 16'hf660;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n18757), .B(\fcw_r_15__N_495[11] ), .C(n18705), 
         .D(n18690), .Z(n16936)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(16[7] 17[28])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h6996;
    FD1S3IX fcw_r_i10 (.D(\fcw_r_15__N_495[11] ), .CK(clk_N_168), .CD(n10972), 
            .Q(fcw_r[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=5, LSE_RCOL=3, LSE_LLINE=146, LSE_RLINE=155 */ ;   // d:/fpga_project/lattice_diamond/piano/dds.v(14[12] 20[6])
    defparam fcw_r_i10.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module sin_rom
//

module sin_rom (\u_count2[24] , \u_count2[23] , \u_count2[22] , \u_count2[21] , 
            \u_count2[20] , \u_count2[19] , \u_count2[18] , \u_count2[17] , 
            \u_count2[16] , \u_count2[15] , \u_count2[14] , clk, \en[1] , 
            GND_net, data_out2, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input \u_count2[24] ;
    input \u_count2[23] ;
    input \u_count2[22] ;
    input \u_count2[21] ;
    input \u_count2[20] ;
    input \u_count2[19] ;
    input \u_count2[18] ;
    input \u_count2[17] ;
    input \u_count2[16] ;
    input \u_count2[15] ;
    input \u_count2[14] ;
    input clk;
    input \en[1] ;
    input GND_net;
    output [11:0]data_out2;
    input VCC_net;
    
    wire clk /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    
    DP8KC sin_rom_0_2_0 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
          .ADA2(\u_count2[14] ), .ADA3(\u_count2[15] ), .ADA4(\u_count2[16] ), 
          .ADA5(\u_count2[17] ), .ADA6(\u_count2[18] ), .ADA7(\u_count2[19] ), 
          .ADA8(\u_count2[20] ), .ADA9(\u_count2[21] ), .ADA10(\u_count2[22] ), 
          .ADA11(\u_count2[23] ), .ADA12(\u_count2[24] ), .CEA(\en[1] ), 
          .OCEA(\en[1] ), .CLKA(clk), .WEA(GND_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(GND_net), 
          .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
          .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
          .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(GND_net), 
          .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
          .RSTB(GND_net), .DOA0(data_out2[8]), .DOA1(data_out2[9]), .DOA2(data_out2[10]), 
          .DOA3(data_out2[11])) /* synthesis MEM_LPC_FILE="sin_rom.lpc", MEM_INIT_FILE="sin_2048.mem", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=38, LSE_RLINE=44 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(38[10] 44[4])
    defparam sin_rom_0_2_0.DATA_WIDTH_A = 4;
    defparam sin_rom_0_2_0.DATA_WIDTH_B = 4;
    defparam sin_rom_0_2_0.REGMODE_A = "OUTREG";
    defparam sin_rom_0_2_0.REGMODE_B = "NOREG";
    defparam sin_rom_0_2_0.CSDECODE_A = "0b000";
    defparam sin_rom_0_2_0.CSDECODE_B = "0b111";
    defparam sin_rom_0_2_0.WRITEMODE_A = "NORMAL";
    defparam sin_rom_0_2_0.WRITEMODE_B = "NORMAL";
    defparam sin_rom_0_2_0.GSR = "ENABLED";
    defparam sin_rom_0_2_0.RESETMODE = "SYNC";
    defparam sin_rom_0_2_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam sin_rom_0_2_0.INIT_DATA = "STATIC";
    defparam sin_rom_0_2_0.INITVAL_00 = "0x176BB176BB176BA154AA154AA154AA154AA152991329913299132991328811088110881108811088";
    defparam sin_rom_0_2_0.INITVAL_01 = "0x1DCEE1DCEE1DADD1BADD1BADD1BADD1BADD1BADD1BACC198CC198CC198CC198CC198CB176BB176BB";
    defparam sin_rom_0_2_0.INITVAL_02 = "0x1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEEE1DCEE1DCEE1DCEE1DCEE1DCEE";
    defparam sin_rom_0_2_0.INITVAL_03 = "0x1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF";
    defparam sin_rom_0_2_0.INITVAL_04 = "0x1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF";
    defparam sin_rom_0_2_0.INITVAL_05 = "0x1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEF1FEFF";
    defparam sin_rom_0_2_0.INITVAL_06 = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_07 = "0x198CC198CC198CC198CC198CC198CC198CC198CC19ADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_08 = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADC198CC198CC198CC198CC198CC198CC198CC198CC198CC";
    defparam sin_rom_0_2_0.INITVAL_09 = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0A = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0B = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0C = "0x198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC19ADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0D = "0x154BB176BB176BB176BB176BB176BB176BB176BB176BB176BB176BB176BB176BB178CC198CC198CC";
    defparam sin_rom_0_2_0.INITVAL_0E = "0x1329913299132991329913299134AA154AA154AA154AA154AA154AA154AA154AA154AA154AA154AA";
    defparam sin_rom_0_2_0.INITVAL_0F = "0x11088110881108811088110881108811088110881108811088110991329913299132991329913299";
    defparam sin_rom_0_2_0.INITVAL_10 = "0x0CC660CC660CC660CC660CC660CE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE78";
    defparam sin_rom_0_2_0.INITVAL_11 = "0x0AA550AA550AA550AA550AA550AA550AA550AA550AA550AA550AA660CC660CC660CC660CC660CC66";
    defparam sin_rom_0_2_0.INITVAL_12 = "0x06633066330664408844088440884408844088440884408844088440884408844088440884408A55";
    defparam sin_rom_0_2_0.INITVAL_13 = "0x04422044330663306633066330663306633066330663306633066330663306633066330663306633";
    defparam sin_rom_0_2_0.INITVAL_14 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_15 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_16 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_17 = "0x06633066330663306633066330663306633066330663306422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_18 = "0x04422044220442204422044220442204422044330663306633066330663306633066330663306633";
    defparam sin_rom_0_2_0.INITVAL_19 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_1A = "0x00000022110221102211022110221102211022110221102211022110221102211022110221102212";
    defparam sin_rom_0_2_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam sin_rom_0_2_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam sin_rom_0_2_0.INITVAL_1D = "0x02211022110221102211022110200000000000000000000000000000000000000000000000000000";
    defparam sin_rom_0_2_0.INITVAL_1E = "0x08844088440663306633066330663306633064220442204422044220442204422044110221102211";
    defparam sin_rom_0_2_0.INITVAL_1F = "0x0EE770EE770EE770EE770EC660CC660CC660CC660CC550AA550AA550AA550AA55088440884408844";
    DP8KC sin_rom_0_0_2 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
          .ADA2(\u_count2[14] ), .ADA3(\u_count2[15] ), .ADA4(\u_count2[16] ), 
          .ADA5(\u_count2[17] ), .ADA6(\u_count2[18] ), .ADA7(\u_count2[19] ), 
          .ADA8(\u_count2[20] ), .ADA9(\u_count2[21] ), .ADA10(\u_count2[22] ), 
          .ADA11(\u_count2[23] ), .ADA12(\u_count2[24] ), .CEA(\en[1] ), 
          .OCEA(\en[1] ), .CLKA(clk), .WEA(GND_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(GND_net), 
          .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
          .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
          .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(GND_net), 
          .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
          .RSTB(GND_net), .DOA0(data_out2[0]), .DOA1(data_out2[1]), .DOA2(data_out2[2]), 
          .DOA3(data_out2[3])) /* synthesis MEM_LPC_FILE="sin_rom.lpc", MEM_INIT_FILE="sin_2048.mem", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=38, LSE_RLINE=44 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(38[10] 44[4])
    defparam sin_rom_0_0_2.DATA_WIDTH_A = 4;
    defparam sin_rom_0_0_2.DATA_WIDTH_B = 4;
    defparam sin_rom_0_0_2.REGMODE_A = "OUTREG";
    defparam sin_rom_0_0_2.REGMODE_B = "NOREG";
    defparam sin_rom_0_0_2.CSDECODE_A = "0b000";
    defparam sin_rom_0_0_2.CSDECODE_B = "0b111";
    defparam sin_rom_0_0_2.WRITEMODE_A = "NORMAL";
    defparam sin_rom_0_0_2.WRITEMODE_B = "NORMAL";
    defparam sin_rom_0_0_2.GSR = "ENABLED";
    defparam sin_rom_0_0_2.RESETMODE = "SYNC";
    defparam sin_rom_0_0_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam sin_rom_0_0_2.INIT_DATA = "STATIC";
    defparam sin_rom_0_0_2.INITVAL_00 = "0x138E106C9B1A0240D2BD1E2350F2AC1C0130AC89178EF004350CE8A178DE0022308A67134BC1BCF0";
    defparam sin_rom_0_0_2.INITVAL_01 = "0x030F61A8B213E6C072F51627D070E413C491C68D04CB0092D10D4E20D4E20B2D008EAE0287A1A036";
    defparam sin_rom_0_0_2.INITVAL_02 = "0x0C60D14C3F190401904016E2E128FA0A0B50145F126E70365E102A41ACF80122A0763B0763B07429";
    defparam sin_rom_0_0_2.INITVAL_03 = "0x08C89178EF024340AC78132AB178CC1BADD1BACC196BA152870CA43040FD194860840E1927405EC9";
    defparam sin_rom_0_0_2.INITVAL_04 = "0x0F6F4118041180411804118F30F6E20D2D008EBE02A8B1C24817C030D2CE0286917C0208E9B1BE13";
    defparam sin_rom_0_0_2.INITVAL_05 = "0x04CAE04EBF06EB0090D10B2E20D6F41181515C27160491A26A1E68C00A9E04CBF090C10B2E20D4F3";
    defparam sin_rom_0_0_2.INITVAL_06 = "0x08C8A1BE240D2BE0266917C140F4DF04C9C1E45819E26138030F4E10B2C008EBF06CAE04CAE04CAE";
    defparam sin_rom_0_0_2.INITVAL_07 = "0x1DEFF1FEFF0000102222066450AC77112AB198DE1E22308A68134CD1E0230AE8A19CF106A7917AF2";
    defparam sin_rom_0_0_2.INITVAL_08 = "0x174980EA430420F1D8BA130760A8330420F1DADC1749910E760CA4406622042100000F1FEFF1FEEE";
    defparam sin_rom_0_0_2.INITVAL_09 = "0x10E650862101EEC174980EC530420F1B8BA12E65084101FACB13076086211FCDB152860A83101EEC";
    defparam sin_rom_0_0_2.INITVAL_0A = "0x1129A154BB198CD1BADD1BCEE1DCEE1DADD1BADC198BB174A9130870EC65088320420F1FCDC17498";
    defparam sin_rom_0_0_2.INITVAL_0B = "0x08C9B1C0350F4CE00657136DF02657114CE002340D09B19AF0046450D09A178DE1E012046450AC77";
    defparam sin_rom_0_0_2.INITVAL_0C = "0x092D10B4E20D4E20D4E20D4E20D4E10B2C008EBF04C9C0067A1A24715A040F4D006C8B1C247138F1";
    defparam sin_rom_0_0_2.INITVAL_0D = "0x11C381C69E072E311C381A68D04ED20F8161605A1E89E070D10D60513C381826A1E68C02AAE06EC0";
    defparam sin_rom_0_0_2.INITVAL_0E = "0x13E5B02EC211C4A00CC20FA391EAB00D8281A69F0B4061627D050E313E4A00AB00D8171847D050D3";
    defparam sin_rom_0_0_2.INITVAL_0F = "0x0D8281CAB10FA391EAB10FC4A00CC211C4A00CC213E5B02ED313E5B02ED313E5B02ED313E5B02ED3";
    defparam sin_rom_0_0_2.INITVAL_10 = "0x072F51627D072F51627D072F51627D072F51627E094061848E094061849F0B6171A69F0B6281C8A0";
    defparam sin_rom_0_0_2.INITVAL_11 = "0x070E313C491E8A00B6061827D050E313E5A00CB10FA381C8A00B6171A69E094061848E092F51627D";
    defparam sin_rom_0_0_2.INITVAL_12 = "0x092D20D6F411A1615E481A47B00AAF070D20F8161605A1E89E072E311A381A48D04ED20FA281A48D";
    defparam sin_rom_0_0_2.INITVAL_13 = "0x0287919E25114D006C9C0066919E3613A040F4E10B2C008EBF04CAE04CAE04CAE04CAE04CBF06EC0";
    defparam sin_rom_0_0_2.INITVAL_14 = "0x134BB19AEE1E012068560F0AB19AE0026450F0AC1BE0208C8917AF106A7917A0208C9B1A0250F4CF";
    defparam sin_rom_0_0_2.INITVAL_15 = "0x0EC540641101EEE1B8CB15499110770CC550A8440663306622044220443306633088450AC660EE89";
    defparam sin_rom_0_0_2.INITVAL_16 = "0x0420F1B8BA10E650641F1DACA13075086101FCCB152760A83101EED174980EC540420F1DACB15288";
    defparam sin_rom_0_0_2.INITVAL_17 = "0x0421102211000001FEEE1DADC196AA132870EC540662101EED1B8BA130760A82101EED196980EC54";
    defparam sin_rom_0_0_2.INITVAL_18 = "0x02657136DF02446112BD1C01308C78156CD1DE12068450CE89134BB19ADE1DEFF000010221102222";
    defparam sin_rom_0_0_2.INITVAL_19 = "0x0D4E20D4E20D4D10B2C008EBF04C9D0087A1C24817C140F4E106C9C1E45715AF20AEAC1C236114CE";
    defparam sin_rom_0_0_2.INITVAL_1A = "0x02CAE04EBF090C10B4E20F60411A1615E37180591C46B1E88C02AAE04EBF070C00B2D10B2E20D4E2";
    defparam sin_rom_0_0_2.INITVAL_1B = "0x1E2350F2CE00457158F208EAD0045819E25116F20B2C006EAE04A9D0288C0088C0088C0088C02A9D";
    defparam sin_rom_0_0_2.INITVAL_1C = "0x082EC12E4201CCA10C43020ED196A910E660AA440863306634088550CE78134BC1BCF104857114CD";
    defparam sin_rom_0_0_2.INITVAL_1D = "0x1CCD51AAD51AAD61CE080343C0DE8216AF905A7116C0B0A0B6038721D25019040190411B46301AA7";
    defparam sin_rom_0_0_2.INITVAL_1E = "0x1A036138F20D2C006EBE04CAE04CAF06EC00B4E311A271847C050D313E5B02ED41427E0B83A030F7";
    defparam sin_rom_0_0_2.INITVAL_1F = "0x024340AC79156CD1DE0206856112AB1BC0104857114BD1E0240CE9B1BE130AEAC1C0350F4DF0487A";
    DP8KC sin_rom_0_1_1 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
          .ADA2(\u_count2[14] ), .ADA3(\u_count2[15] ), .ADA4(\u_count2[16] ), 
          .ADA5(\u_count2[17] ), .ADA6(\u_count2[18] ), .ADA7(\u_count2[19] ), 
          .ADA8(\u_count2[20] ), .ADA9(\u_count2[21] ), .ADA10(\u_count2[22] ), 
          .ADA11(\u_count2[23] ), .ADA12(\u_count2[24] ), .CEA(\en[1] ), 
          .OCEA(\en[1] ), .CLKA(clk), .WEA(GND_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(GND_net), 
          .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
          .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
          .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(GND_net), 
          .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
          .RSTB(GND_net), .DOA0(data_out2[4]), .DOA1(data_out2[5]), .DOA2(data_out2[6]), 
          .DOA3(data_out2[7])) /* synthesis MEM_LPC_FILE="sin_rom.lpc", MEM_INIT_FILE="sin_2048.mem", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=38, LSE_RLINE=44 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(38[10] 44[4])
    defparam sin_rom_0_1_1.DATA_WIDTH_A = 4;
    defparam sin_rom_0_1_1.DATA_WIDTH_B = 4;
    defparam sin_rom_0_1_1.REGMODE_A = "OUTREG";
    defparam sin_rom_0_1_1.REGMODE_B = "NOREG";
    defparam sin_rom_0_1_1.CSDECODE_A = "0b000";
    defparam sin_rom_0_1_1.CSDECODE_B = "0b111";
    defparam sin_rom_0_1_1.WRITEMODE_A = "NORMAL";
    defparam sin_rom_0_1_1.WRITEMODE_B = "NORMAL";
    defparam sin_rom_0_1_1.GSR = "ENABLED";
    defparam sin_rom_0_1_1.RESETMODE = "SYNC";
    defparam sin_rom_0_1_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam sin_rom_0_1_1.INIT_DATA = "STATIC";
    defparam sin_rom_0_1_1.INITVAL_00 = "0x10E660A8320220F1DACB154980EC540662101EED196A9130760A832020FE1DACB152870CA4304200";
    defparam sin_rom_0_1_1.INITVAL_01 = "0x0A8330441101EFE1DACC176A9130770CA5406621020FF1DACC1749910E660A8330420F1FCDC176A9";
    defparam sin_rom_0_1_1.INITVAL_02 = "0x198CB176BA154AA13299110870EE660CC550A8430662204210000FF1DCDD1B8CB174A9130870EC65";
    defparam sin_rom_0_1_1.INITVAL_03 = "0x1DCEE1DCEE1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEEE1DCEE1DCED1BADD1B8CC";
    defparam sin_rom_0_1_1.INITVAL_04 = "0x022120443306644088550AA560CC670EE781108813299134AA154BB176BB198CC198DD1BADD1BAEE";
    defparam sin_rom_0_1_1.INITVAL_05 = "0x00000022110442306634088450AA560CC770EE8811299134AA156BB198CC1BADD1DCEF1FEF000001";
    defparam sin_rom_0_1_1.INITVAL_06 = "0x0663306644088440AA550AA660CC660EE770F08811099132AA154AB176BC198CC1BADD1DCEE1FEFF";
    defparam sin_rom_0_1_1.INITVAL_07 = "0x1DCEE1DCEE1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1E00000000000000021102211022120442204423";
    defparam sin_rom_0_1_1.INITVAL_08 = "0x0221102211022100000000000000000000F1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFE1DCEE1DCEE";
    defparam sin_rom_0_1_1.INITVAL_09 = "0x0CC660CC660CA550AA550AA550AA5408844088440884406633066330663304422044220442204211";
    defparam sin_rom_0_1_1.INITVAL_0A = "0x0EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE760CC660CC66";
    defparam sin_rom_0_1_1.INITVAL_0B = "0x022110242204422066330663308844088440AA550AA550AA560CC660CC660CC660CE770EE770EE77";
    defparam sin_rom_0_1_1.INITVAL_0C = "0x06634088450AA560CC670EE78110891329A154AA176BB198CC19ADD1BAEE1DCEF1FEFF1E00000001";
    defparam sin_rom_0_1_1.INITVAL_0D = "0x1FE0000211044230664408A550CC670EE8811299134AA176BC198DD1BAEE1DEFF1E0000221104423";
    defparam sin_rom_0_1_1.INITVAL_0E = "0x11099154AB176CC1BADE1DCFF1E0010222204633088550AC660EE7811099154AB176CC19ADD1DCEF";
    defparam sin_rom_0_1_1.INITVAL_0F = "0x00011024230664408A560CC7711089132AA176BC198DD1DCEF1FE000221204433088450AA660EE78";
    defparam sin_rom_0_1_1.INITVAL_10 = "0x11089134AA176BC19ADD1DCEF1E0000221204633088550AC660EE8811299154BB178CC1BAEE1DEF0";
    defparam sin_rom_0_1_1.INITVAL_11 = "0x0221204433068450AA660CE7711089132AA176BC198DD1BCEF1FE000021104433068440AA560CE77";
    defparam sin_rom_0_1_1.INITVAL_12 = "0x1BADE1DCEF1FE00000110242206633088450AA660CE770F0881329A154BB178CC1BADE1DCFF1E000";
    defparam sin_rom_0_1_1.INITVAL_13 = "0x1FEFF1FE000000102211044220443306644088450AA560CC660EE771108813299154AA176BB198CD";
    defparam sin_rom_0_1_1.INITVAL_14 = "0x11088110881129913299132991329A154AA154AA154BB176BB176BC198CC198DD1BADD1BCEE1DCEE";
    defparam sin_rom_0_1_1.INITVAL_15 = "0x13299132991308811088110881108811088110881108811088110881108811088110881108811088";
    defparam sin_rom_0_1_1.INITVAL_16 = "0x1DCED1BADD1BADD1BADC198CC198CC198CC176BB176BB176BB174AA154AA154AA154A91329913299";
    defparam sin_rom_0_1_1.INITVAL_17 = "0x02211022110221100000000000000000000000000000001EFF1FEFF1FEFF1FEFF1FCEE1DCEE1DCEE";
    defparam sin_rom_0_1_1.INITVAL_18 = "0x1BADD1BADD1DCEE1DCEE1DEFF1FEFF1FEFF1FE000000000000000000000000000022110221102211";
    defparam sin_rom_0_1_1.INITVAL_19 = "0x00001022120442306634088440AA550CC660CE770EE881108913299134AA154AB176BB178CC198CC";
    defparam sin_rom_0_1_1.INITVAL_1A = "0x1FEFF00000022120442306644088550AA660CE770F08811299154AA176BB198CD1BADE1DCEF1FEF0";
    defparam sin_rom_0_1_1.INITVAL_1B = "0x02422044220663306634088440AA550AA660CC670EE781108813299154AA176BB198CC1BADD1DCEE";
    defparam sin_rom_0_1_1.INITVAL_1C = "0x06622044220421102211022000000000000000000000000000000000000000000000010221102211";
    defparam sin_rom_0_1_1.INITVAL_1D = "0x132880EE660AA44066320421001EFF1DCDD1B8CC176BA15499130880EE770CC660AA550884408633";
    defparam sin_rom_0_1_1.INITVAL_1E = "0x0AA43042001FCDD196A9130760CA430641101EEE1B8CB1549810E660A84306411000FE1DADC196AA";
    defparam sin_rom_0_1_1.INITVAL_1F = "0x1FCDC174980EC540642101EED196A910E760A832020FE1BACB152870CA54064101FEED196A913076";
    
endmodule
//
// Verilog Description of module sin_rom_U12
//

module sin_rom_U12 (\u_count1[24] , \u_count1[23] , \u_count1[22] , \u_count1[21] , 
            \u_count1[20] , \u_count1[19] , \u_count1[18] , \u_count1[17] , 
            \u_count1[16] , \u_count1[15] , \u_count1[14] , clk, \en[0] , 
            GND_net, data_out1, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input \u_count1[24] ;
    input \u_count1[23] ;
    input \u_count1[22] ;
    input \u_count1[21] ;
    input \u_count1[20] ;
    input \u_count1[19] ;
    input \u_count1[18] ;
    input \u_count1[17] ;
    input \u_count1[16] ;
    input \u_count1[15] ;
    input \u_count1[14] ;
    input clk;
    input \en[0] ;
    input GND_net;
    output [11:0]data_out1;
    input VCC_net;
    
    wire clk /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    
    DP8KC sin_rom_0_2_0 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
          .ADA2(\u_count1[14] ), .ADA3(\u_count1[15] ), .ADA4(\u_count1[16] ), 
          .ADA5(\u_count1[17] ), .ADA6(\u_count1[18] ), .ADA7(\u_count1[19] ), 
          .ADA8(\u_count1[20] ), .ADA9(\u_count1[21] ), .ADA10(\u_count1[22] ), 
          .ADA11(\u_count1[23] ), .ADA12(\u_count1[24] ), .CEA(\en[0] ), 
          .OCEA(\en[0] ), .CLKA(clk), .WEA(GND_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(GND_net), 
          .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
          .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
          .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(GND_net), 
          .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
          .RSTB(GND_net), .DOA0(data_out1[8]), .DOA1(data_out1[9]), .DOA2(data_out1[10]), 
          .DOA3(data_out1[11])) /* synthesis MEM_LPC_FILE="sin_rom.lpc", MEM_INIT_FILE="sin_2048.mem", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=31, LSE_RLINE=37 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(31[10] 37[4])
    defparam sin_rom_0_2_0.DATA_WIDTH_A = 4;
    defparam sin_rom_0_2_0.DATA_WIDTH_B = 4;
    defparam sin_rom_0_2_0.REGMODE_A = "OUTREG";
    defparam sin_rom_0_2_0.REGMODE_B = "NOREG";
    defparam sin_rom_0_2_0.CSDECODE_A = "0b000";
    defparam sin_rom_0_2_0.CSDECODE_B = "0b111";
    defparam sin_rom_0_2_0.WRITEMODE_A = "NORMAL";
    defparam sin_rom_0_2_0.WRITEMODE_B = "NORMAL";
    defparam sin_rom_0_2_0.GSR = "ENABLED";
    defparam sin_rom_0_2_0.RESETMODE = "SYNC";
    defparam sin_rom_0_2_0.ASYNC_RESET_RELEASE = "SYNC";
    defparam sin_rom_0_2_0.INIT_DATA = "STATIC";
    defparam sin_rom_0_2_0.INITVAL_00 = "0x176BB176BB176BA154AA154AA154AA154AA152991329913299132991328811088110881108811088";
    defparam sin_rom_0_2_0.INITVAL_01 = "0x1DCEE1DCEE1DADD1BADD1BADD1BADD1BADD1BADD1BACC198CC198CC198CC198CC198CB176BB176BB";
    defparam sin_rom_0_2_0.INITVAL_02 = "0x1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEEE1DCEE1DCEE1DCEE1DCEE1DCEE";
    defparam sin_rom_0_2_0.INITVAL_03 = "0x1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF";
    defparam sin_rom_0_2_0.INITVAL_04 = "0x1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF";
    defparam sin_rom_0_2_0.INITVAL_05 = "0x1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEE1DCEF1FEFF";
    defparam sin_rom_0_2_0.INITVAL_06 = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_07 = "0x198CC198CC198CC198CC198CC198CC198CC198CC19ADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_08 = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADC198CC198CC198CC198CC198CC198CC198CC198CC198CC";
    defparam sin_rom_0_2_0.INITVAL_09 = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0A = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0B = "0x1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0C = "0x198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC198CC19ADD1BADD";
    defparam sin_rom_0_2_0.INITVAL_0D = "0x154BB176BB176BB176BB176BB176BB176BB176BB176BB176BB176BB176BB176BB178CC198CC198CC";
    defparam sin_rom_0_2_0.INITVAL_0E = "0x1329913299132991329913299134AA154AA154AA154AA154AA154AA154AA154AA154AA154AA154AA";
    defparam sin_rom_0_2_0.INITVAL_0F = "0x11088110881108811088110881108811088110881108811088110991329913299132991329913299";
    defparam sin_rom_0_2_0.INITVAL_10 = "0x0CC660CC660CC660CC660CC660CE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE78";
    defparam sin_rom_0_2_0.INITVAL_11 = "0x0AA550AA550AA550AA550AA550AA550AA550AA550AA550AA550AA660CC660CC660CC660CC660CC66";
    defparam sin_rom_0_2_0.INITVAL_12 = "0x06633066330664408844088440884408844088440884408844088440884408844088440884408A55";
    defparam sin_rom_0_2_0.INITVAL_13 = "0x04422044330663306633066330663306633066330663306633066330663306633066330663306633";
    defparam sin_rom_0_2_0.INITVAL_14 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_15 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_16 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_17 = "0x06633066330663306633066330663306633066330663306422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_18 = "0x04422044220442204422044220442204422044330663306633066330663306633066330663306633";
    defparam sin_rom_0_2_0.INITVAL_19 = "0x04422044220442204422044220442204422044220442204422044220442204422044220442204422";
    defparam sin_rom_0_2_0.INITVAL_1A = "0x00000022110221102211022110221102211022110221102211022110221102211022110221102212";
    defparam sin_rom_0_2_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam sin_rom_0_2_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam sin_rom_0_2_0.INITVAL_1D = "0x02211022110221102211022110200000000000000000000000000000000000000000000000000000";
    defparam sin_rom_0_2_0.INITVAL_1E = "0x08844088440663306633066330663306633064220442204422044220442204422044110221102211";
    defparam sin_rom_0_2_0.INITVAL_1F = "0x0EE770EE770EE770EE770EC660CC660CC660CC660CC550AA550AA550AA550AA55088440884408844";
    DP8KC sin_rom_0_1_1 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
          .ADA2(\u_count1[14] ), .ADA3(\u_count1[15] ), .ADA4(\u_count1[16] ), 
          .ADA5(\u_count1[17] ), .ADA6(\u_count1[18] ), .ADA7(\u_count1[19] ), 
          .ADA8(\u_count1[20] ), .ADA9(\u_count1[21] ), .ADA10(\u_count1[22] ), 
          .ADA11(\u_count1[23] ), .ADA12(\u_count1[24] ), .CEA(\en[0] ), 
          .OCEA(\en[0] ), .CLKA(clk), .WEA(GND_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(GND_net), 
          .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
          .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
          .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(GND_net), 
          .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
          .RSTB(GND_net), .DOA0(data_out1[4]), .DOA1(data_out1[5]), .DOA2(data_out1[6]), 
          .DOA3(data_out1[7])) /* synthesis MEM_LPC_FILE="sin_rom.lpc", MEM_INIT_FILE="sin_2048.mem", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=31, LSE_RLINE=37 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(31[10] 37[4])
    defparam sin_rom_0_1_1.DATA_WIDTH_A = 4;
    defparam sin_rom_0_1_1.DATA_WIDTH_B = 4;
    defparam sin_rom_0_1_1.REGMODE_A = "OUTREG";
    defparam sin_rom_0_1_1.REGMODE_B = "NOREG";
    defparam sin_rom_0_1_1.CSDECODE_A = "0b000";
    defparam sin_rom_0_1_1.CSDECODE_B = "0b111";
    defparam sin_rom_0_1_1.WRITEMODE_A = "NORMAL";
    defparam sin_rom_0_1_1.WRITEMODE_B = "NORMAL";
    defparam sin_rom_0_1_1.GSR = "ENABLED";
    defparam sin_rom_0_1_1.RESETMODE = "SYNC";
    defparam sin_rom_0_1_1.ASYNC_RESET_RELEASE = "SYNC";
    defparam sin_rom_0_1_1.INIT_DATA = "STATIC";
    defparam sin_rom_0_1_1.INITVAL_00 = "0x10E660A8320220F1DACB154980EC540662101EED196A9130760A832020FE1DACB152870CA4304200";
    defparam sin_rom_0_1_1.INITVAL_01 = "0x0A8330441101EFE1DACC176A9130770CA5406621020FF1DACC1749910E660A8330420F1FCDC176A9";
    defparam sin_rom_0_1_1.INITVAL_02 = "0x198CB176BA154AA13299110870EE660CC550A8430662204210000FF1DCDD1B8CB174A9130870EC65";
    defparam sin_rom_0_1_1.INITVAL_03 = "0x1DCEE1DCEE1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEEE1DCEE1DCED1BADD1B8CC";
    defparam sin_rom_0_1_1.INITVAL_04 = "0x022120443306644088550AA560CC670EE781108813299134AA154BB176BB198CC198DD1BADD1BAEE";
    defparam sin_rom_0_1_1.INITVAL_05 = "0x00000022110442306634088450AA560CC770EE8811299134AA156BB198CC1BADD1DCEF1FEF000001";
    defparam sin_rom_0_1_1.INITVAL_06 = "0x0663306644088440AA550AA660CC660EE770F08811099132AA154AB176BC198CC1BADD1DCEE1FEFF";
    defparam sin_rom_0_1_1.INITVAL_07 = "0x1DCEE1DCEE1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1E00000000000000021102211022120442204423";
    defparam sin_rom_0_1_1.INITVAL_08 = "0x0221102211022100000000000000000000F1FEFF1FEFF1FEFF1FEFF1FEFF1FEFF1FEFE1DCEE1DCEE";
    defparam sin_rom_0_1_1.INITVAL_09 = "0x0CC660CC660CA550AA550AA550AA5408844088440884406633066330663304422044220442204211";
    defparam sin_rom_0_1_1.INITVAL_0A = "0x0EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE770EE760CC660CC66";
    defparam sin_rom_0_1_1.INITVAL_0B = "0x022110242204422066330663308844088440AA550AA550AA560CC660CC660CC660CE770EE770EE77";
    defparam sin_rom_0_1_1.INITVAL_0C = "0x06634088450AA560CC670EE78110891329A154AA176BB198CC19ADD1BAEE1DCEF1FEFF1E00000001";
    defparam sin_rom_0_1_1.INITVAL_0D = "0x1FE0000211044230664408A550CC670EE8811299134AA176BC198DD1BAEE1DEFF1E0000221104423";
    defparam sin_rom_0_1_1.INITVAL_0E = "0x11099154AB176CC1BADE1DCFF1E0010222204633088550AC660EE7811099154AB176CC19ADD1DCEF";
    defparam sin_rom_0_1_1.INITVAL_0F = "0x00011024230664408A560CC7711089132AA176BC198DD1DCEF1FE000221204433088450AA660EE78";
    defparam sin_rom_0_1_1.INITVAL_10 = "0x11089134AA176BC19ADD1DCEF1E0000221204633088550AC660EE8811299154BB178CC1BAEE1DEF0";
    defparam sin_rom_0_1_1.INITVAL_11 = "0x0221204433068450AA660CE7711089132AA176BC198DD1BCEF1FE000021104433068440AA560CE77";
    defparam sin_rom_0_1_1.INITVAL_12 = "0x1BADE1DCEF1FE00000110242206633088450AA660CE770F0881329A154BB178CC1BADE1DCFF1E000";
    defparam sin_rom_0_1_1.INITVAL_13 = "0x1FEFF1FE000000102211044220443306644088450AA560CC660EE771108813299154AA176BB198CD";
    defparam sin_rom_0_1_1.INITVAL_14 = "0x11088110881129913299132991329A154AA154AA154BB176BB176BC198CC198DD1BADD1BCEE1DCEE";
    defparam sin_rom_0_1_1.INITVAL_15 = "0x13299132991308811088110881108811088110881108811088110881108811088110881108811088";
    defparam sin_rom_0_1_1.INITVAL_16 = "0x1DCED1BADD1BADD1BADC198CC198CC198CC176BB176BB176BB174AA154AA154AA154A91329913299";
    defparam sin_rom_0_1_1.INITVAL_17 = "0x02211022110221100000000000000000000000000000001EFF1FEFF1FEFF1FEFF1FCEE1DCEE1DCEE";
    defparam sin_rom_0_1_1.INITVAL_18 = "0x1BADD1BADD1DCEE1DCEE1DEFF1FEFF1FEFF1FE000000000000000000000000000022110221102211";
    defparam sin_rom_0_1_1.INITVAL_19 = "0x00001022120442306634088440AA550CC660CE770EE881108913299134AA154AB176BB178CC198CC";
    defparam sin_rom_0_1_1.INITVAL_1A = "0x1FEFF00000022120442306644088550AA660CE770F08811299154AA176BB198CD1BADE1DCEF1FEF0";
    defparam sin_rom_0_1_1.INITVAL_1B = "0x02422044220663306634088440AA550AA660CC670EE781108813299154AA176BB198CC1BADD1DCEE";
    defparam sin_rom_0_1_1.INITVAL_1C = "0x06622044220421102211022000000000000000000000000000000000000000000000010221102211";
    defparam sin_rom_0_1_1.INITVAL_1D = "0x132880EE660AA44066320421001EFF1DCDD1B8CC176BA15499130880EE770CC660AA550884408633";
    defparam sin_rom_0_1_1.INITVAL_1E = "0x0AA43042001FCDD196A9130760CA430641101EEE1B8CB1549810E660A84306411000FE1DADC196AA";
    defparam sin_rom_0_1_1.INITVAL_1F = "0x1FCDC174980EC540642101EED196A910E760A832020FE1BACB152870CA54064101FEED196A913076";
    DP8KC sin_rom_0_0_2 (.DIA0(GND_net), .DIA1(GND_net), .DIA2(GND_net), 
          .DIA3(GND_net), .DIA4(GND_net), .DIA5(GND_net), .DIA6(GND_net), 
          .DIA7(GND_net), .DIA8(GND_net), .ADA0(GND_net), .ADA1(GND_net), 
          .ADA2(\u_count1[14] ), .ADA3(\u_count1[15] ), .ADA4(\u_count1[16] ), 
          .ADA5(\u_count1[17] ), .ADA6(\u_count1[18] ), .ADA7(\u_count1[19] ), 
          .ADA8(\u_count1[20] ), .ADA9(\u_count1[21] ), .ADA10(\u_count1[22] ), 
          .ADA11(\u_count1[23] ), .ADA12(\u_count1[24] ), .CEA(\en[0] ), 
          .OCEA(\en[0] ), .CLKA(clk), .WEA(GND_net), .CSA0(GND_net), 
          .CSA1(GND_net), .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), 
          .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), 
          .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), 
          .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(GND_net), 
          .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), .ADB7(GND_net), 
          .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), .ADB11(GND_net), 
          .ADB12(GND_net), .CEB(VCC_net), .OCEB(VCC_net), .CLKB(GND_net), 
          .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
          .RSTB(GND_net), .DOA0(data_out1[0]), .DOA1(data_out1[1]), .DOA2(data_out1[2]), 
          .DOA3(data_out1[3])) /* synthesis MEM_LPC_FILE="sin_rom.lpc", MEM_INIT_FILE="sin_2048.mem", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=31, LSE_RLINE=37 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(31[10] 37[4])
    defparam sin_rom_0_0_2.DATA_WIDTH_A = 4;
    defparam sin_rom_0_0_2.DATA_WIDTH_B = 4;
    defparam sin_rom_0_0_2.REGMODE_A = "OUTREG";
    defparam sin_rom_0_0_2.REGMODE_B = "NOREG";
    defparam sin_rom_0_0_2.CSDECODE_A = "0b000";
    defparam sin_rom_0_0_2.CSDECODE_B = "0b111";
    defparam sin_rom_0_0_2.WRITEMODE_A = "NORMAL";
    defparam sin_rom_0_0_2.WRITEMODE_B = "NORMAL";
    defparam sin_rom_0_0_2.GSR = "ENABLED";
    defparam sin_rom_0_0_2.RESETMODE = "SYNC";
    defparam sin_rom_0_0_2.ASYNC_RESET_RELEASE = "SYNC";
    defparam sin_rom_0_0_2.INIT_DATA = "STATIC";
    defparam sin_rom_0_0_2.INITVAL_00 = "0x138E106C9B1A0240D2BD1E2350F2AC1C0130AC89178EF004350CE8A178DE0022308A67134BC1BCF0";
    defparam sin_rom_0_0_2.INITVAL_01 = "0x030F61A8B213E6C072F51627D070E413C491C68D04CB0092D10D4E20D4E20B2D008EAE0287A1A036";
    defparam sin_rom_0_0_2.INITVAL_02 = "0x0C60D14C3F190401904016E2E128FA0A0B50145F126E70365E102A41ACF80122A0763B0763B07429";
    defparam sin_rom_0_0_2.INITVAL_03 = "0x08C89178EF024340AC78132AB178CC1BADD1BACC196BA152870CA43040FD194860840E1927405EC9";
    defparam sin_rom_0_0_2.INITVAL_04 = "0x0F6F4118041180411804118F30F6E20D2D008EBE02A8B1C24817C030D2CE0286917C0208E9B1BE13";
    defparam sin_rom_0_0_2.INITVAL_05 = "0x04CAE04EBF06EB0090D10B2E20D6F41181515C27160491A26A1E68C00A9E04CBF090C10B2E20D4F3";
    defparam sin_rom_0_0_2.INITVAL_06 = "0x08C8A1BE240D2BE0266917C140F4DF04C9C1E45819E26138030F4E10B2C008EBF06CAE04CAE04CAE";
    defparam sin_rom_0_0_2.INITVAL_07 = "0x1DEFF1FEFF0000102222066450AC77112AB198DE1E22308A68134CD1E0230AE8A19CF106A7917AF2";
    defparam sin_rom_0_0_2.INITVAL_08 = "0x174980EA430420F1D8BA130760A8330420F1DADC1749910E760CA4406622042100000F1FEFF1FEEE";
    defparam sin_rom_0_0_2.INITVAL_09 = "0x10E650862101EEC174980EC530420F1B8BA12E65084101FACB13076086211FCDB152860A83101EEC";
    defparam sin_rom_0_0_2.INITVAL_0A = "0x1129A154BB198CD1BADD1BCEE1DCEE1DADD1BADC198BB174A9130870EC65088320420F1FCDC17498";
    defparam sin_rom_0_0_2.INITVAL_0B = "0x08C9B1C0350F4CE00657136DF02657114CE002340D09B19AF0046450D09A178DE1E012046450AC77";
    defparam sin_rom_0_0_2.INITVAL_0C = "0x092D10B4E20D4E20D4E20D4E20D4E10B2C008EBF04C9C0067A1A24715A040F4D006C8B1C247138F1";
    defparam sin_rom_0_0_2.INITVAL_0D = "0x11C381C69E072E311C381A68D04ED20F8161605A1E89E070D10D60513C381826A1E68C02AAE06EC0";
    defparam sin_rom_0_0_2.INITVAL_0E = "0x13E5B02EC211C4A00CC20FA391EAB00D8281A69F0B4061627D050E313E4A00AB00D8171847D050D3";
    defparam sin_rom_0_0_2.INITVAL_0F = "0x0D8281CAB10FA391EAB10FC4A00CC211C4A00CC213E5B02ED313E5B02ED313E5B02ED313E5B02ED3";
    defparam sin_rom_0_0_2.INITVAL_10 = "0x072F51627D072F51627D072F51627D072F51627E094061848E094061849F0B6171A69F0B6281C8A0";
    defparam sin_rom_0_0_2.INITVAL_11 = "0x070E313C491E8A00B6061827D050E313E5A00CB10FA381C8A00B6171A69E094061848E092F51627D";
    defparam sin_rom_0_0_2.INITVAL_12 = "0x092D20D6F411A1615E481A47B00AAF070D20F8161605A1E89E072E311A381A48D04ED20FA281A48D";
    defparam sin_rom_0_0_2.INITVAL_13 = "0x0287919E25114D006C9C0066919E3613A040F4E10B2C008EBF04CAE04CAE04CAE04CAE04CBF06EC0";
    defparam sin_rom_0_0_2.INITVAL_14 = "0x134BB19AEE1E012068560F0AB19AE0026450F0AC1BE0208C8917AF106A7917A0208C9B1A0250F4CF";
    defparam sin_rom_0_0_2.INITVAL_15 = "0x0EC540641101EEE1B8CB15499110770CC550A8440663306622044220443306633088450AC660EE89";
    defparam sin_rom_0_0_2.INITVAL_16 = "0x0420F1B8BA10E650641F1DACA13075086101FCCB152760A83101EED174980EC540420F1DACB15288";
    defparam sin_rom_0_0_2.INITVAL_17 = "0x0421102211000001FEEE1DADC196AA132870EC540662101EED1B8BA130760A82101EED196980EC54";
    defparam sin_rom_0_0_2.INITVAL_18 = "0x02657136DF02446112BD1C01308C78156CD1DE12068450CE89134BB19ADE1DEFF000010221102222";
    defparam sin_rom_0_0_2.INITVAL_19 = "0x0D4E20D4E20D4D10B2C008EBF04C9D0087A1C24817C140F4E106C9C1E45715AF20AEAC1C236114CE";
    defparam sin_rom_0_0_2.INITVAL_1A = "0x02CAE04EBF090C10B4E20F60411A1615E37180591C46B1E88C02AAE04EBF070C00B2D10B2E20D4E2";
    defparam sin_rom_0_0_2.INITVAL_1B = "0x1E2350F2CE00457158F208EAD0045819E25116F20B2C006EAE04A9D0288C0088C0088C0088C02A9D";
    defparam sin_rom_0_0_2.INITVAL_1C = "0x082EC12E4201CCA10C43020ED196A910E660AA440863306634088550CE78134BC1BCF104857114CD";
    defparam sin_rom_0_0_2.INITVAL_1D = "0x1CCD51AAD51AAD61CE080343C0DE8216AF905A7116C0B0A0B6038721D25019040190411B46301AA7";
    defparam sin_rom_0_0_2.INITVAL_1E = "0x1A036138F20D2C006EBE04CAE04CAF06EC00B4E311A271847C050D313E5B02ED41427E0B83A030F7";
    defparam sin_rom_0_0_2.INITVAL_1F = "0x024340AC79156CD1DE0206856112AB1BC0104857114BD1E0240CE9B1BE130AEAC1C0350F4DF0487A";
    
endmodule
//
// Verilog Description of module key
//

module key (clk_N_168, key_state_flag, key_state_c, key_state_value, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output key_state_flag;
    input key_state_c;
    output key_state_value;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18788, n10399, key_flag_N_639, key_reg, n15528;
    wire [31:0]n9;
    
    wire n15527, n15526, n15525, n15524, n15523, n15522, n15521, 
        n15520, n15519, n15518, n15517, n15516, n15515, n15514, 
        n15513, n10264, clk_N_168_enable_505, clk_N_168_enable_493;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n55, n60, n49, n50, n48, n39_adj_829, n58, n52, n40_adj_830, 
        n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10399), .CK(clk_N_168), .CD(n18788), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(key_state_flag)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_state_c), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_state_c), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(key_state_value)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15528), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15527), .COUT(n15528), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15526), .COUT(n15527), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15525), .COUT(n15526), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15524), .COUT(n15525), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15523), .COUT(n15524), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15522), .COUT(n15523), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15521), .COUT(n15522), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15520), .COUT(n15521), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15519), .COUT(n15520), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15518), .COUT(n15519), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15517), .COUT(n15518), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15516), .COUT(n15517), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15515), .COUT(n15516), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15514), .COUT(n15515), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15513), .COUT(n15514), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15513), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i5555_2_lut_rep_442 (.A(delay_cnt[0]), .B(n10264), .Z(clk_N_168_enable_505)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5555_2_lut_rep_442.init = 16'heeee;
    LUT4 i5556_2_lut_3_lut (.A(delay_cnt[0]), .B(n10264), .C(n9[0]), .Z(n10399)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5556_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_493), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_505), .CD(n18788), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=172, LSE_RLINE=178 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    LUT4 key_reg_I_0_2_lut_rep_606 (.A(key_reg), .B(key_state_c), .Z(n18788)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_606.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_state_c), .C(n10264), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_493)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i7531_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[19]), 
         .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7531_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7530_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[18]), 
         .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7530_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7529_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[17]), 
         .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7529_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7528_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[16]), 
         .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7528_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7527_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[14]), 
         .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7527_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7526_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7526_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7525_2_lut_3_lut (.A(key_reg), .B(key_state_c), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7525_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10264)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_829), .B(n58), .C(n52), .D(n40_adj_830), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_829)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_830)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12327_2_lut (.A(delay_cnt[0]), .B(n10264), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12327_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module buzzer
//

module buzzer (CNT, GND_net, CNT_17__N_703, clk_N_168, stat, \yinjie_box_2__N_394[0] , 
            \yinjie_box_2__N_394[1] , n77, n9292, n19846, \data_out2[0] , 
            \data_out1[0] , n28, yinjie, pwm_out1_c, \PWM_in_12__N_452[12] , 
            \PWM_in_12__N_452[11] , \PWM_in_12__N_452[10] , \rom2[0] , 
            n18850, \PWM_in_12__N_452[9] , n97, n18725, n18707, n18706, 
            n18709, n18721, n18616, \cycle_17__N_740[4] , n17110, 
            n18755, n18708, n18736, n18684, n7, \cycle_17__N_740[13] , 
            \PWM_in_12__N_452[8] , n407, \cycle_17__N_740[11] , n18722, 
            n18763, \cycle_17__N_740[14] , n415, \cycle_17__N_740[3] , 
            \note[0] , n18737, n18807, n18697, n18757, n18784, n18785, 
            \fcw_r_15__N_495[8] , \PWM_in_12__N_452[7] , n18690, \fcw_r_15__N_495[6] , 
            n8146, n8147, \fcw_r_15__N_495[10] , \fcw_r_15__N_495[5] , 
            n18717, n10972, \fcw_r_15__N_495[11] , \fcw_r_15__N_495[9] , 
            n18620, n18668, n16876, \cycle_17__N_740[1] , \note[1] , 
            n18808, n12983, \PWM_in_12__N_452[6] , \PWM_in_12__N_452[5] , 
            n406, \cycle_17__N_740[12] , clk_N_168_enable_507, \cycle_17__N_663[2] , 
            clk_N_168_enable_512, \cycle_17__N_663[7] , \cycle_17__N_663[10] , 
            clk_N_168_enable_518, \cycle_17__N_663[17] , \cycle_17__N_740[9] , 
            n18769, \PWM_in_12__N_452[4] , n19_adj_4, n22_adj_5, n18772, 
            n14_adj_6, n3, n3_adj_7, n18735, n16828, n18754, n262, 
            \PWM_in_12__N_452[3] , n7_adj_8, \cycle_17__N_740[16] , \PWM_in_12__N_452[2] , 
            n18720, n18815, n18651, \PWM_in_12__N_452[1] , n18803, 
            n18761, n18768, n18771, n18619, clk__inv, n410, n18623, 
            \key_value[0] , \key_value[10] , n269, n16959, n26_adj_9, 
            n9757, \cycle_17__N_740[10] , n18308, n18307, \key_value[12] , 
            \key_value[5] , \key_value[1] , \key_value[8] , \key_value[7] , 
            \key_value[6] , \key_value[2] , \key_value[11] , \key_value[3] , 
            \key_value[4] , \key_value[9] , n3830, n18679, n436, n18676, 
            \rom1_4__N_338[0] , n351, n414, n31, n18682, n16888, 
            n18610, n247, n331, \rom2[1] , \key_flag[2] , \key_flag[1] , 
            n18734, rst_n_c, key_pa_c, n19839, n18680, n9, n9654, 
            n10160, n344, n18696, n18606, n18612, n16920, n10337, 
            n18649, n18685, n18652, n16909) /* synthesis syn_module_defined=1 */ ;
    output [17:0]CNT;
    input GND_net;
    output [18:0]CNT_17__N_703;
    input clk_N_168;
    input stat;
    input \yinjie_box_2__N_394[0] ;
    input \yinjie_box_2__N_394[1] ;
    output [17:0]n77;
    output n9292;
    input n19846;
    input \data_out2[0] ;
    input \data_out1[0] ;
    output [12:0]n28;
    input [2:0]yinjie;
    output pwm_out1_c;
    input \PWM_in_12__N_452[12] ;
    input \PWM_in_12__N_452[11] ;
    input \PWM_in_12__N_452[10] ;
    input \rom2[0] ;
    output n18850;
    input \PWM_in_12__N_452[9] ;
    input [17:0]n97;
    input n18725;
    input n18707;
    input n18706;
    input n18709;
    input n18721;
    input n18616;
    input \cycle_17__N_740[4] ;
    input n17110;
    input n18755;
    input n18708;
    input n18736;
    input n18684;
    input n7;
    input \cycle_17__N_740[13] ;
    input \PWM_in_12__N_452[8] ;
    input n407;
    input \cycle_17__N_740[11] ;
    input n18722;
    input n18763;
    input \cycle_17__N_740[14] ;
    input n415;
    input \cycle_17__N_740[3] ;
    input \note[0] ;
    input n18737;
    input n18807;
    input n18697;
    output n18757;
    input n18784;
    input n18785;
    output \fcw_r_15__N_495[8] ;
    input \PWM_in_12__N_452[7] ;
    output n18690;
    output \fcw_r_15__N_495[6] ;
    output n8146;
    output n8147;
    output \fcw_r_15__N_495[10] ;
    output \fcw_r_15__N_495[5] ;
    output n18717;
    output n10972;
    output \fcw_r_15__N_495[11] ;
    output \fcw_r_15__N_495[9] ;
    input n18620;
    input n18668;
    output n16876;
    input \cycle_17__N_740[1] ;
    input \note[1] ;
    input n18808;
    input n12983;
    input \PWM_in_12__N_452[6] ;
    input \PWM_in_12__N_452[5] ;
    input n406;
    input \cycle_17__N_740[12] ;
    input clk_N_168_enable_507;
    input \cycle_17__N_663[2] ;
    input clk_N_168_enable_512;
    input \cycle_17__N_663[7] ;
    input \cycle_17__N_663[10] ;
    input clk_N_168_enable_518;
    input \cycle_17__N_663[17] ;
    input \cycle_17__N_740[9] ;
    output n18769;
    input \PWM_in_12__N_452[4] ;
    input n19_adj_4;
    input n22_adj_5;
    output n18772;
    output n14_adj_6;
    input n3;
    input n3_adj_7;
    input n18735;
    output n16828;
    input n18754;
    output n262;
    input \PWM_in_12__N_452[3] ;
    input n7_adj_8;
    input \cycle_17__N_740[16] ;
    input \PWM_in_12__N_452[2] ;
    input n18720;
    input n18815;
    output n18651;
    input \PWM_in_12__N_452[1] ;
    output n18803;
    input n18761;
    input n18768;
    input n18771;
    output n18619;
    input clk__inv;
    input n410;
    input n18623;
    input \key_value[0] ;
    input \key_value[10] ;
    input n269;
    input n16959;
    output n26_adj_9;
    input n9757;
    output \cycle_17__N_740[10] ;
    input n18308;
    input n18307;
    input \key_value[12] ;
    input \key_value[5] ;
    input \key_value[1] ;
    input \key_value[8] ;
    input \key_value[7] ;
    input \key_value[6] ;
    input \key_value[2] ;
    input \key_value[11] ;
    input \key_value[3] ;
    input \key_value[4] ;
    input \key_value[9] ;
    input n3830;
    input n18679;
    input n436;
    input n18676;
    output \rom1_4__N_338[0] ;
    input n351;
    output n414;
    output n31;
    input n18682;
    input n16888;
    input n18610;
    input n247;
    output n331;
    input \rom2[1] ;
    input \key_flag[2] ;
    input \key_flag[1] ;
    output n18734;
    input rst_n_c;
    input key_pa_c;
    output n19839;
    input n18680;
    input n9;
    input n9654;
    input n10160;
    output n344;
    input n18696;
    input n18606;
    input n18612;
    input n16920;
    input n10337;
    input n18649;
    input n18685;
    input n18652;
    input n16909;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire clk__inv /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire [17:0]cycle;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(13[12:17])
    
    wire n12, n30, n15307, n15308, clk_N_168_enable_15;
    wire [17:0]cycle_17__N_663;
    wire [2:0]yinjie_box;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(15[11:21])
    
    wire n15782, n15781, n15780, n15779, n15778, n15777, n15776, 
        n15775, n15774, PWM, n15306, n18848, n18849, n18740, n17088, 
        pwm_out1_N_122, n18739, n14_adj_801, n18741, n26_adj_802, 
        n18742, n18743, n17066, n18, n18744, n20, n14161, n24, 
        n32, n17091, n34, n7_c, n17413, n17071, n18745, n4, 
        n18748, n4_adj_805, n28_c, n17081, n18738, n17097, n10, 
        n18749, n18751, n17052, n8, n18752, n16_adj_806, n17028, 
        n18640, n6, n6_adj_807, n18650, n7_adj_808, n15951, PWM_N_764;
    wire [17:0]cycle_17__N_740;
    
    wire clk_N_168_enable_511, n7_adj_809, clk_N_168_enable_508, clk_N_168_enable_509, 
        clk_N_168_enable_510, clk_N_168_enable_513, clk_N_168_enable_514, 
        clk_N_168_enable_515, clk_N_168_enable_516, clk_N_168_enable_517, 
        clk_N_168_enable_520, clk_N_168_enable_522, n7_adj_811;
    wire [17:0]n400;
    
    wire n17069, n17411, n17050, n15314, n15313, n18648, n17037, 
        n11, n14162, n22_adj_818, n7_adj_819, n15312, n15311, n15310, 
        n24_adj_820, n20_adj_821, n22_adj_823, n16_adj_824, n15309, 
        n29, n17345, n30_adj_825, n31_adj_826, n28_adj_827, n18617, 
        n8_adj_828;
    
    LUT4 CNT_17__I_0_91_i30_3_lut_3_lut (.A(CNT[16]), .B(cycle[17]), .C(n12), 
         .Z(n30)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i30_3_lut_3_lut.init = 16'hd4d4;
    CCU2D sub_6_add_2_5 (.A0(cycle[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cycle[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15307), 
          .COUT(n15308), .S0(CNT_17__N_703[3]), .S1(CNT_17__N_703[4]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_5.INIT0 = 16'h5555;
    defparam sub_6_add_2_5.INIT1 = 16'h5555;
    defparam sub_6_add_2_5.INJECT1_0 = "NO";
    defparam sub_6_add_2_5.INJECT1_1 = "NO";
    FD1P3AX cycle_i0 (.D(cycle_17__N_663[0]), .SP(clk_N_168_enable_15), 
            .CK(clk_N_168), .Q(cycle[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i0.GSR = "DISABLED";
    FD1P3AY yinjie_box_i0 (.D(\yinjie_box_2__N_394[0] ), .SP(stat), .CK(clk_N_168), 
            .Q(yinjie_box[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(93[8] 105[5])
    defparam yinjie_box_i0.GSR = "DISABLED";
    FD1P3AX yinjie_box_i1 (.D(\yinjie_box_2__N_394[1] ), .SP(stat), .CK(clk_N_168), 
            .Q(yinjie_box[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(93[8] 105[5])
    defparam yinjie_box_i1.GSR = "DISABLED";
    CCU2D CNT_2225_add_4_19 (.A0(CNT[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15782), .S0(n77[17]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_19.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_19.INIT1 = 16'h0000;
    defparam CNT_2225_add_4_19.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_19.INJECT1_1 = "NO";
    LUT4 i7345_3_lut_4_lut (.A(n9292), .B(n19846), .C(\data_out2[0] ), 
         .D(\data_out1[0] ), .Z(n28[0])) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7345_3_lut_4_lut.init = 16'h0dd0;
    CCU2D CNT_2225_add_4_17 (.A0(CNT[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15781), .COUT(n15782), .S0(n77[15]), .S1(n77[16]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_17.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_17.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_17.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_17.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_15 (.A0(CNT[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15780), .COUT(n15781), .S0(n77[13]), .S1(n77[14]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_15.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_15.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_15.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_15.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_13 (.A0(CNT[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15779), .COUT(n15780), .S0(n77[11]), .S1(n77[12]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_13.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_13.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_13.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_13.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_11 (.A0(CNT[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15778), .COUT(n15779), .S0(n77[9]), .S1(n77[10]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_11.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_11.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_11.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_11.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_9 (.A0(CNT[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(CNT[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15777), 
          .COUT(n15778), .S0(n77[7]), .S1(n77[8]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_9.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_9.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_9.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_9.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_7 (.A0(CNT[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(CNT[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15776), 
          .COUT(n15777), .S0(n77[5]), .S1(n77[6]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_7.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_7.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_7.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_7.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_5 (.A0(CNT[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(CNT[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15775), 
          .COUT(n15776), .S0(n77[3]), .S1(n77[4]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_5.INIT0 = 16'hfaaa;
    defparam CNT_2225_add_4_5.INIT1 = 16'hfaaa;
    defparam CNT_2225_add_4_5.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_5.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_3 (.A0(CNT[1]), .B0(n19846), .C0(yinjie_box[1]), 
          .D0(yinjie[1]), .A1(yinjie[2]), .B1(n19846), .C1(CNT[2]), 
          .D1(GND_net), .CIN(n15774), .COUT(n15775), .S0(n77[1]), .S1(n77[2]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_3.INIT0 = 16'h596a;
    defparam CNT_2225_add_4_3.INIT1 = 16'hd2d2;
    defparam CNT_2225_add_4_3.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_3.INJECT1_1 = "NO";
    CCU2D CNT_2225_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(CNT[0]), .B1(n19846), .C1(yinjie_box[0]), 
          .D1(yinjie[0]), .COUT(n15774), .S1(n77[0]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225_add_4_1.INIT0 = 16'hF000;
    defparam CNT_2225_add_4_1.INIT1 = 16'h596a;
    defparam CNT_2225_add_4_1.INJECT1_0 = "NO";
    defparam CNT_2225_add_4_1.INJECT1_1 = "NO";
    LUT4 i7314_2_lut_3_lut (.A(n9292), .B(n19846), .C(PWM), .Z(pwm_out1_c)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7314_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7761_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[12] ), 
         .Z(n28[12])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7761_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7760_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[11] ), 
         .Z(n28[11])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7760_2_lut_3_lut.init = 16'hd0d0;
    CCU2D sub_6_add_2_3 (.A0(cycle[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cycle[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15306), 
          .COUT(n15307), .S0(CNT_17__N_703[1]), .S1(CNT_17__N_703[2]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_3.INIT0 = 16'h5555;
    defparam sub_6_add_2_3.INIT1 = 16'h5555;
    defparam sub_6_add_2_3.INJECT1_0 = "NO";
    defparam sub_6_add_2_3.INJECT1_1 = "NO";
    LUT4 i7759_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[10] ), 
         .Z(n28[10])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7759_2_lut_3_lut.init = 16'hd0d0;
    PFUMX i12622 (.BLUT(n18848), .ALUT(n18849), .C0(\rom2[0] ), .Z(n18850));
    LUT4 i7758_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[9] ), 
         .Z(n28[9])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7758_2_lut_3_lut.init = 16'hd0d0;
    LUT4 CNT_17__I_0_91_i29_2_lut_rep_558 (.A(CNT[14]), .B(cycle[15]), .Z(n18740)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i29_2_lut_rep_558.init = 16'h6666;
    LUT4 i11797_2_lut_3_lut_4_lut (.A(CNT[14]), .B(cycle[15]), .C(cycle[14]), 
         .D(CNT[13]), .Z(n17088)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11797_2_lut_3_lut_4_lut.init = 16'h9009;
    FD1S3DX CNT_2225__i0 (.D(n97[0]), .CK(clk_N_168), .CD(pwm_out1_N_122), 
            .Q(CNT[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i0.GSR = "DISABLED";
    LUT4 CNT_17__I_0_91_i27_2_lut_rep_557 (.A(CNT[13]), .B(cycle[14]), .Z(n18739)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i27_2_lut_rep_557.init = 16'h6666;
    LUT4 CNT_17__I_0_91_i14_3_lut_3_lut (.A(CNT[14]), .B(cycle[15]), .C(cycle[14]), 
         .Z(n14_adj_801)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i14_3_lut_3_lut.init = 16'hd4d4;
    LUT4 CNT_17__I_0_91_i31_2_lut_rep_559 (.A(CNT[15]), .B(cycle[16]), .Z(n18741)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i31_2_lut_rep_559.init = 16'h6666;
    LUT4 CNT_17__I_0_91_i26_3_lut_3_lut (.A(CNT[15]), .B(cycle[16]), .C(n14_adj_801), 
         .Z(n26_adj_802)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i26_3_lut_3_lut.init = 16'hd4d4;
    LUT4 CNT_17__I_0_91_i21_2_lut_rep_560 (.A(CNT[10]), .B(cycle[11]), .Z(n18742)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i21_2_lut_rep_560.init = 16'h6666;
    LUT4 CNT_17__I_0_91_i23_2_lut_rep_561 (.A(CNT[11]), .B(cycle[12]), .Z(n18743)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i23_2_lut_rep_561.init = 16'h6666;
    LUT4 i11775_2_lut_3_lut_4_lut (.A(CNT[11]), .B(cycle[12]), .C(cycle[11]), 
         .D(CNT[10]), .Z(n17066)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11775_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 CNT_17__I_0_91_i18_3_lut_3_lut (.A(CNT[11]), .B(cycle[12]), .C(cycle[11]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 CNT_17__I_0_91_i25_2_lut_rep_562 (.A(CNT[12]), .B(cycle[13]), .Z(n18744)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i25_2_lut_rep_562.init = 16'h6666;
    LUT4 CNT_17__I_0_91_i20_3_lut_3_lut (.A(CNT[12]), .B(cycle[13]), .C(n18), 
         .Z(n20)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i8_3_lut_4_lut (.A(n18725), .B(n18707), .C(n18706), .D(n18709), 
         .Z(n14161)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(47[4] 48[25])
    defparam i8_3_lut_4_lut.init = 16'h0001;
    LUT4 i2_3_lut_4_lut (.A(n18725), .B(n18707), .C(n18721), .D(n18616), 
         .Z(clk_N_168_enable_15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(47[4] 48[25])
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    L6MUX21 CNT_17__I_0_91_i34 (.D0(n24), .D1(n32), .SD(n17091), .Z(n34)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    PFUMX mux_57_i5 (.BLUT(n7_c), .ALUT(\cycle_17__N_740[4] ), .C0(n17110), 
          .Z(cycle_17__N_663[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 i12354_2_lut_3_lut (.A(CNT[12]), .B(cycle[13]), .C(n17413), .Z(n17071)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12354_2_lut_3_lut.init = 16'hf6f6;
    LUT4 CNT_17__I_0_91_i9_2_lut_rep_563 (.A(CNT[4]), .B(cycle[5]), .Z(n18745)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i9_2_lut_rep_563.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n18755), .B(n18708), .C(n18736), .D(n18684), 
         .Z(n4)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(63[4] 64[24])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hefee;
    PFUMX mux_57_i14 (.BLUT(n7), .ALUT(\cycle_17__N_740[13] ), .C0(n17110), 
          .Z(cycle_17__N_663[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 i7757_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[8] ), 
         .Z(n28[8])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7757_2_lut_3_lut.init = 16'hd0d0;
    LUT4 CNT_17__I_0_91_i13_2_lut_rep_566 (.A(CNT[6]), .B(cycle[7]), .Z(n18748)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i13_2_lut_rep_566.init = 16'h6666;
    LUT4 i12182_4_lut_4_lut (.A(n18741), .B(n17088), .C(n26_adj_802), 
         .D(n4_adj_805), .Z(n28_c)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12182_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i12348_4_lut_4_lut (.A(n18741), .B(n17081), .C(n18740), .D(n18738), 
         .Z(n17097)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12348_4_lut_4_lut.init = 16'hff04;
    LUT4 CNT_17__I_0_91_i10_3_lut_3_lut (.A(CNT[6]), .B(cycle[7]), .C(cycle[6]), 
         .Z(n10)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 CNT_17__I_0_91_i15_2_lut_rep_567 (.A(CNT[7]), .B(cycle[8]), .Z(n18749)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i15_2_lut_rep_567.init = 16'h6666;
    LUT4 CNT_17__I_0_91_i12_3_lut_3_lut (.A(CNT[7]), .B(cycle[8]), .C(n10), 
         .Z(n12)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 CNT_17__I_0_91_i17_2_lut_rep_569 (.A(CNT[8]), .B(cycle[9]), .Z(n18751)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i17_2_lut_rep_569.init = 16'h6666;
    LUT4 i11761_2_lut_3_lut_4_lut (.A(CNT[8]), .B(cycle[9]), .C(cycle[5]), 
         .D(CNT[4]), .Z(n17052)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11761_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 CNT_17__I_0_91_i8_3_lut_3_lut (.A(CNT[8]), .B(cycle[9]), .C(cycle[5]), 
         .Z(n8)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 CNT_17__I_0_91_i19_2_lut_rep_570 (.A(CNT[9]), .B(cycle[10]), .Z(n18752)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i19_2_lut_rep_570.init = 16'h6666;
    LUT4 CNT_17__I_0_91_i16_3_lut_3_lut (.A(CNT[9]), .B(cycle[10]), .C(n8), 
         .Z(n16_adj_806)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i16_3_lut_3_lut.init = 16'hd4d4;
    PFUMX mux_57_i12 (.BLUT(n407), .ALUT(\cycle_17__N_740[11] ), .C0(n19846), 
          .Z(cycle_17__N_663[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 i11737_3_lut_4_lut (.A(CNT[3]), .B(cycle[4]), .C(cycle[3]), .D(CNT[2]), 
         .Z(n17028)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11737_3_lut_4_lut.init = 16'h9009;
    LUT4 i1_2_lut_rep_458_3_lut_4_lut (.A(n18721), .B(n18725), .C(n18736), 
         .D(n18722), .Z(n18640)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_458_3_lut_4_lut.init = 16'hfffe;
    LUT4 CNT_17__I_0_91_i6_3_lut_3_lut (.A(CNT[3]), .B(cycle[4]), .C(cycle[3]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_3_lut_4_lut_adj_17 (.A(n18721), .B(n18725), .C(n19846), 
         .D(n18763), .Z(n6_adj_807)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_17.init = 16'hfffe;
    LUT4 i1_2_lut_rep_468_3_lut_4_lut (.A(n18725), .B(n18722), .C(n18721), 
         .D(n19846), .Z(n18650)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(45[4] 46[25])
    defparam i1_2_lut_rep_468_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_57_i15 (.BLUT(n7_adj_808), .ALUT(\cycle_17__N_740[14] ), .C0(n17110), 
          .Z(cycle_17__N_663[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    FD1S3JX PWM_89 (.D(PWM_N_764), .CK(clk_N_168), .PD(n15951), .Q(PWM)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(108[8] 115[4])
    defparam PWM_89.GSR = "DISABLED";
    PFUMX mux_57_i4 (.BLUT(n415), .ALUT(\cycle_17__N_740[3] ), .C0(n19846), 
          .Z(cycle_17__N_663[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 i2_4_lut_4_lut (.A(\note[0] ), .B(n18737), .C(n18807), .D(n18697), 
         .Z(cycle_17__N_740[8])) /* synthesis lut_function=(A (C (D))+!A !((C+!(D))+!B)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i2_4_lut_4_lut.init = 16'ha400;
    LUT4 i7373_2_lut_rep_575 (.A(yinjie[2]), .B(n19846), .Z(n18757)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i7373_2_lut_rep_575.init = 16'h2222;
    LUT4 i3039_2_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), 
         .C(n18784), .D(n18785), .Z(\fcw_r_15__N_495[8] )) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (D)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i3039_2_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hdd20;
    LUT4 i7756_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[7] ), 
         .Z(n28[7])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7756_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i4128_2_lut_rep_508_4_lut (.A(yinjie[2]), .B(n19846), .C(n18784), 
         .D(n18785), .Z(n18690)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i4128_2_lut_rep_508_4_lut.init = 16'hd200;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), 
         .C(n18784), .D(n18785), .Z(\fcw_r_15__N_495[6] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A ((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h20d2;
    LUT4 i4006_3_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), .C(n18785), 
         .D(n18784), .Z(n8146)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i4006_3_lut_3_lut_4_lut.init = 16'h2ff0;
    LUT4 i3998_2_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), .C(n18785), 
         .D(n18784), .Z(n8147)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i3998_2_lut_3_lut_4_lut.init = 16'hd2f0;
    LUT4 i3188_2_lut_rep_464_3_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), 
         .C(n18784), .D(n18785), .Z(\fcw_r_15__N_495[10] )) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i3188_2_lut_rep_464_3_lut_3_lut_4_lut.init = 16'h0222;
    LUT4 i4126_2_lut_3_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), .C(n18784), 
         .D(n18785), .Z(\fcw_r_15__N_495[5] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (C (D)+!C !(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i4126_2_lut_3_lut_3_lut_4_lut.init = 16'h2df0;
    LUT4 i10322_2_lut_rep_535_4_lut (.A(yinjie[2]), .B(n19846), .C(n18785), 
         .D(n18784), .Z(n18717)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i10322_2_lut_rep_535_4_lut.init = 16'h2d22;
    LUT4 i6114_1_lut_2_lut (.A(yinjie[2]), .B(n19846), .Z(n10972)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i6114_1_lut_2_lut.init = 16'hdddd;
    LUT4 CNT_17__I_0_91_i4_4_lut (.A(cycle[1]), .B(cycle[2]), .C(CNT[1]), 
         .D(CNT[0]), .Z(n4_adj_805)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A ((C)+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i4_4_lut.init = 16'h0c8e;
    LUT4 i3784_2_lut_3_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), .C(n18784), 
         .D(n18785), .Z(\fcw_r_15__N_495[11] )) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i3784_2_lut_3_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i3047_2_lut_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(yinjie[2]), .B(n19846), 
         .C(n18784), .D(n18785), .Z(\fcw_r_15__N_495[9] )) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i3047_2_lut_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hd2f0;
    LUT4 i1_2_lut_4_lut (.A(n18620), .B(n18763), .C(n18668), .D(n16876), 
         .Z(clk_N_168_enable_511)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(65[4] 66[24])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    PFUMX mux_57_i2 (.BLUT(n7_adj_809), .ALUT(\cycle_17__N_740[1] ), .C0(n17110), 
          .Z(cycle_17__N_663[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 CNT_17__I_0_91_i33_2_lut_rep_556 (.A(CNT[16]), .B(cycle[17]), .Z(n18738)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i33_2_lut_rep_556.init = 16'h6666;
    LUT4 mux_63_Mux_6_i15_4_lut_4_lut (.A(\note[1] ), .B(n18808), .C(n18807), 
         .D(n12983), .Z(cycle_17__N_740[6])) /* synthesis lut_function=(!(A (C)+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_6_i15_4_lut_4_lut.init = 16'h4f4a;
    LUT4 i7755_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[6] ), 
         .Z(n28[6])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7755_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i7754_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[5] ), 
         .Z(n28[5])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7754_2_lut_3_lut.init = 16'hd0d0;
    PFUMX mux_57_i13 (.BLUT(n406), .ALUT(\cycle_17__N_740[12] ), .C0(n19846), 
          .Z(cycle_17__N_663[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    FD1P3AX cycle_i1 (.D(cycle_17__N_663[1]), .SP(clk_N_168_enable_508), 
            .CK(clk_N_168), .Q(cycle[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i1.GSR = "DISABLED";
    FD1P3AX cycle_i2 (.D(\cycle_17__N_663[2] ), .SP(clk_N_168_enable_507), 
            .CK(clk_N_168), .Q(cycle[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i2.GSR = "DISABLED";
    FD1P3AX cycle_i3 (.D(cycle_17__N_663[3]), .SP(clk_N_168_enable_508), 
            .CK(clk_N_168), .Q(cycle[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i3.GSR = "DISABLED";
    FD1P3AX cycle_i4 (.D(cycle_17__N_663[4]), .SP(clk_N_168_enable_509), 
            .CK(clk_N_168), .Q(cycle[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i4.GSR = "DISABLED";
    FD1P3AX cycle_i5 (.D(cycle_17__N_663[5]), .SP(clk_N_168_enable_510), 
            .CK(clk_N_168), .Q(cycle[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i5.GSR = "DISABLED";
    FD1P3AX cycle_i6 (.D(cycle_17__N_663[6]), .SP(clk_N_168_enable_511), 
            .CK(clk_N_168), .Q(cycle[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i6.GSR = "DISABLED";
    FD1P3AX cycle_i7 (.D(\cycle_17__N_663[7] ), .SP(clk_N_168_enable_512), 
            .CK(clk_N_168), .Q(cycle[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i7.GSR = "DISABLED";
    FD1P3AX cycle_i8 (.D(cycle_17__N_663[8]), .SP(clk_N_168_enable_513), 
            .CK(clk_N_168), .Q(cycle[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i8.GSR = "DISABLED";
    FD1P3AX cycle_i9 (.D(cycle_17__N_663[9]), .SP(clk_N_168_enable_514), 
            .CK(clk_N_168), .Q(cycle[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i9.GSR = "DISABLED";
    FD1P3AX cycle_i10 (.D(\cycle_17__N_663[10] ), .SP(clk_N_168_enable_515), 
            .CK(clk_N_168), .Q(cycle[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i10.GSR = "DISABLED";
    FD1P3AX cycle_i11 (.D(cycle_17__N_663[11]), .SP(clk_N_168_enable_516), 
            .CK(clk_N_168), .Q(cycle[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i11.GSR = "DISABLED";
    FD1P3AX cycle_i12 (.D(cycle_17__N_663[12]), .SP(clk_N_168_enable_517), 
            .CK(clk_N_168), .Q(cycle[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i12.GSR = "DISABLED";
    FD1P3AX cycle_i13 (.D(cycle_17__N_663[13]), .SP(clk_N_168_enable_518), 
            .CK(clk_N_168), .Q(cycle[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i13.GSR = "DISABLED";
    FD1P3AX cycle_i14 (.D(cycle_17__N_663[14]), .SP(clk_N_168_enable_520), 
            .CK(clk_N_168), .Q(cycle[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i14.GSR = "DISABLED";
    FD1P3AX cycle_i15 (.D(cycle_17__N_663[15]), .SP(clk_N_168_enable_520), 
            .CK(clk_N_168), .Q(cycle[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i15.GSR = "DISABLED";
    FD1P3AX cycle_i16 (.D(cycle_17__N_663[16]), .SP(clk_N_168_enable_522), 
            .CK(clk_N_168), .Q(cycle[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i16.GSR = "DISABLED";
    FD1P3AX cycle_i17 (.D(\cycle_17__N_663[17] ), .SP(clk_N_168_enable_522), 
            .CK(clk_N_168), .Q(cycle[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(39[7] 90[4])
    defparam cycle_i17.GSR = "DISABLED";
    PFUMX mux_57_i10 (.BLUT(n7_adj_811), .ALUT(\cycle_17__N_740[9] ), .C0(n17110), 
          .Z(cycle_17__N_663[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    PFUMX mux_57_i7 (.BLUT(n400[6]), .ALUT(cycle_17__N_740[6]), .C0(n19846), 
          .Z(cycle_17__N_663[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 i2985_2_lut_rep_587 (.A(\note[0] ), .B(\note[1] ), .Z(n18769)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i2985_2_lut_rep_587.init = 16'h6666;
    LUT4 i12351_4_lut (.A(n18741), .B(n18740), .C(n18739), .D(n17069), 
         .Z(n17411)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12351_4_lut.init = 16'hfffe;
    LUT4 i7753_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[4] ), 
         .Z(n28[4])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7753_2_lut_3_lut.init = 16'hd0d0;
    PFUMX CNT_17__I_0_91_i32 (.BLUT(n28_c), .ALUT(n30), .C0(n17097), .Z(n32)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    PFUMX i38 (.BLUT(n19_adj_4), .ALUT(n22_adj_5), .C0(n17110), .Z(cycle_17__N_663[15]));
    LUT4 i12260_2_lut_rep_590 (.A(\note[0] ), .B(\note[1] ), .Z(n18772)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i12260_2_lut_rep_590.init = 16'h9999;
    LUT4 i7812_2_lut_3_lut (.A(\note[0] ), .B(\note[1] ), .C(n18808), 
         .Z(n14_adj_6)) /* synthesis lut_function=(A (B (C))+!A !(B+!(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i7812_2_lut_3_lut.init = 16'h9090;
    LUT4 mux_63_Mux_14_i7_3_lut_3_lut_4_lut (.A(\note[0] ), .B(\note[1] ), 
         .C(n3), .D(n18808), .Z(n7_adj_808)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_14_i7_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_63_Mux_9_i7_3_lut_3_lut_4_lut (.A(\note[0] ), .B(\note[1] ), 
         .C(n3_adj_7), .D(n18808), .Z(n7_adj_811)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_9_i7_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i11778_4_lut (.A(n18744), .B(n18743), .C(n18742), .D(n17050), 
         .Z(n17069)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11778_4_lut.init = 16'h0100;
    CCU2D sub_6_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cycle[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n15306), 
          .S1(CNT_17__N_703[0]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_1.INIT0 = 16'hF000;
    defparam sub_6_add_2_1.INIT1 = 16'h5555;
    defparam sub_6_add_2_1.INJECT1_0 = "NO";
    defparam sub_6_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_6_add_2_19 (.A0(cycle[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15314), .S0(CNT_17__N_703[17]), .S1(CNT_17__N_703[18]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_19.INIT0 = 16'h5555;
    defparam sub_6_add_2_19.INIT1 = 16'hffff;
    defparam sub_6_add_2_19.INJECT1_0 = "NO";
    defparam sub_6_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_6_add_2_17 (.A0(cycle[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15313), .COUT(n15314), .S0(CNT_17__N_703[15]), 
          .S1(CNT_17__N_703[16]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_17.INIT0 = 16'h5555;
    defparam sub_6_add_2_17.INIT1 = 16'h5555;
    defparam sub_6_add_2_17.INJECT1_0 = "NO";
    defparam sub_6_add_2_17.INJECT1_1 = "NO";
    LUT4 mux_63_Mux_0_i15_4_lut (.A(\note[0] ), .B(n18808), .C(n18807), 
         .D(\note[1] ), .Z(cycle_17__N_740[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_0_i15_4_lut.init = 16'hc2c8;
    LUT4 i1_3_lut_4_lut (.A(n18736), .B(n18722), .C(n18725), .D(n18735), 
         .Z(n16828)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(47[4] 48[25])
    defparam i1_3_lut_4_lut.init = 16'h00ef;
    LUT4 i6074_2_lut_3_lut_4_lut (.A(n18736), .B(n18722), .C(n18735), 
         .D(n18754), .Z(n262)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(47[4] 48[25])
    defparam i6074_2_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_2_lut_rep_466_3_lut_4_lut (.A(n18736), .B(n18722), .C(n18725), 
         .D(n18721), .Z(n18648)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(47[4] 48[25])
    defparam i1_2_lut_rep_466_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12352_2_lut_3_lut (.A(CNT[16]), .B(cycle[17]), .C(n17411), .Z(n17091)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12352_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7752_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[3] ), 
         .Z(n28[3])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7752_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i11759_4_lut (.A(n18752), .B(n18751), .C(n18749), .D(n17037), 
         .Z(n17050)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11759_4_lut.init = 16'h1011;
    LUT4 i11746_4_lut (.A(n18748), .B(n11), .C(n18745), .D(n17028), 
         .Z(n17037)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11746_4_lut.init = 16'h1011;
    PFUMX mux_57_i17 (.BLUT(n7_adj_8), .ALUT(\cycle_17__N_740[16] ), .C0(n17110), 
          .Z(cycle_17__N_663[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 mux_63_Mux_1_i7_3_lut_3_lut_4_lut (.A(\note[0] ), .B(\note[1] ), 
         .C(n3_adj_7), .D(n18808), .Z(n7_adj_809)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_1_i7_3_lut_3_lut_4_lut.init = 16'hf022;
    LUT4 i7751_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[2] ), 
         .Z(n28[2])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7751_2_lut_3_lut.init = 16'hd0d0;
    PFUMX i9369 (.BLUT(n14161), .ALUT(cycle_17__N_740[0]), .C0(n19846), 
          .Z(n14162));
    LUT4 i1_2_lut_rep_469_3_lut_4_lut (.A(n18720), .B(n18815), .C(n18735), 
         .D(n18754), .Z(n18651)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(63[4] 64[24])
    defparam i1_2_lut_rep_469_3_lut_4_lut.init = 16'hfffe;
    PFUMX CNT_17__I_0_91_i24 (.BLUT(n16_adj_806), .ALUT(n22_adj_818), .C0(n17071), 
          .Z(n24)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 i7750_2_lut_3_lut (.A(n9292), .B(n19846), .C(\PWM_in_12__N_452[1] ), 
         .Z(n28[1])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(117[18:63])
    defparam i7750_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i12335_2_lut_rep_621 (.A(\note[0] ), .B(\note[1] ), .Z(n18803)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i12335_2_lut_rep_621.init = 16'h1111;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\note[0] ), .B(\note[1] ), .C(n18808), 
         .Z(n7_adj_819)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i1_2_lut_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_437_2_lut_3_lut_3_lut_4_lut (.A(n18761), .B(n18763), 
         .C(n18768), .D(n18771), .Z(n18619)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_437_2_lut_3_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12163_4_lut_4_lut (.A(n18744), .B(n17066), .C(n20), .D(n6), 
         .Z(n22_adj_818)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12163_4_lut_4_lut.init = 16'hf4b0;
    FD1S3DX CNT_2225__i1 (.D(n97[1]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i1.GSR = "DISABLED";
    FD1S3DX CNT_2225__i2 (.D(n97[2]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i2.GSR = "DISABLED";
    FD1S3DX CNT_2225__i3 (.D(n97[3]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i3.GSR = "DISABLED";
    FD1S3DX CNT_2225__i4 (.D(n97[4]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i4.GSR = "DISABLED";
    FD1S3DX CNT_2225__i5 (.D(n97[5]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i5.GSR = "DISABLED";
    FD1S3DX CNT_2225__i6 (.D(n97[6]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i6.GSR = "DISABLED";
    FD1S3DX CNT_2225__i7 (.D(n97[7]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i7.GSR = "DISABLED";
    FD1S3DX CNT_2225__i8 (.D(n97[8]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i8.GSR = "DISABLED";
    FD1S3DX CNT_2225__i9 (.D(n97[9]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i9.GSR = "DISABLED";
    FD1S3DX CNT_2225__i10 (.D(n97[10]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i10.GSR = "DISABLED";
    FD1S3DX CNT_2225__i11 (.D(n97[11]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i11.GSR = "DISABLED";
    FD1S3DX CNT_2225__i12 (.D(n97[12]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i12.GSR = "DISABLED";
    FD1S3DX CNT_2225__i13 (.D(n97[13]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i13.GSR = "DISABLED";
    FD1S3DX CNT_2225__i14 (.D(n97[14]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i14.GSR = "DISABLED";
    FD1S3DX CNT_2225__i15 (.D(n97[15]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i15.GSR = "DISABLED";
    FD1S3DX CNT_2225__i16 (.D(n97[16]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i16.GSR = "DISABLED";
    FD1S3DX CNT_2225__i17 (.D(n97[17]), .CK(clk__inv), .CD(pwm_out1_N_122), 
            .Q(CNT[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam CNT_2225__i17.GSR = "DISABLED";
    CCU2D sub_6_add_2_15 (.A0(cycle[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15312), .COUT(n15313), .S0(CNT_17__N_703[13]), 
          .S1(CNT_17__N_703[14]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_15.INIT0 = 16'h5555;
    defparam sub_6_add_2_15.INIT1 = 16'h5555;
    defparam sub_6_add_2_15.INJECT1_0 = "NO";
    defparam sub_6_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_6_add_2_13 (.A0(cycle[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15311), .COUT(n15312), .S0(CNT_17__N_703[11]), 
          .S1(CNT_17__N_703[12]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_13.INIT0 = 16'h5555;
    defparam sub_6_add_2_13.INIT1 = 16'h5555;
    defparam sub_6_add_2_13.INJECT1_0 = "NO";
    defparam sub_6_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_6_add_2_11 (.A0(cycle[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cycle[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15310), .COUT(n15311), .S0(CNT_17__N_703[9]), .S1(CNT_17__N_703[10]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_11.INIT0 = 16'h5555;
    defparam sub_6_add_2_11.INIT1 = 16'h5555;
    defparam sub_6_add_2_11.INJECT1_0 = "NO";
    defparam sub_6_add_2_11.INJECT1_1 = "NO";
    PFUMX mux_57_i9 (.BLUT(n410), .ALUT(cycle_17__N_740[8]), .C0(n19846), 
          .Z(cycle_17__N_663[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=182, LSE_RLINE=191 */ ;
    LUT4 mux_63_Mux_4_i7_3_lut_3_lut_3_lut (.A(\note[0] ), .B(\note[1] ), 
         .C(n18808), .Z(n7_c)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_4_i7_3_lut_3_lut_3_lut.init = 16'hc2c2;
    LUT4 CNT_17__I_0_91_i11_2_lut (.A(CNT[5]), .B(cycle[6]), .Z(n11)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam CNT_17__I_0_91_i11_2_lut.init = 16'h6666;
    LUT4 i1_4_lut (.A(n14162), .B(n18709), .C(n18623), .D(n19846), .Z(cycle_17__N_663[0])) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'haaba;
    LUT4 i12_4_lut (.A(\key_value[0] ), .B(n24_adj_820), .C(n20_adj_821), 
         .D(\key_value[10] ), .Z(n9292)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12_4_lut.init = 16'h8000;
    LUT4 i12353_4_lut (.A(n18743), .B(n18742), .C(n18752), .D(n17052), 
         .Z(n17413)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i12353_4_lut.init = 16'hefee;
    LUT4 i1_4_lut_adj_18 (.A(n18709), .B(n269), .C(n16959), .D(n18720), 
         .Z(n26_adj_9)) /* synthesis lut_function=(A+!(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_18.init = 16'hafae;
    LUT4 i7546_4_lut (.A(n18706), .B(n18763), .C(n18620), .D(n4), .Z(n400[6])) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(65[4] 66[24])
    defparam i7546_4_lut.init = 16'hcfce;
    LUT4 mux_63_Mux_10_i15_4_lut (.A(n7_adj_819), .B(\note[0] ), .C(n18807), 
         .D(n9757), .Z(\cycle_17__N_740[10] )) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam mux_63_Mux_10_i15_4_lut.init = 16'h0a3a;
    PFUMX i12480 (.BLUT(n18308), .ALUT(n18307), .C0(n19846), .Z(cycle_17__N_663[5]));
    LUT4 i11_4_lut (.A(\key_value[12] ), .B(n22_adj_823), .C(n16_adj_824), 
         .D(\key_value[5] ), .Z(n24_adj_820)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11_4_lut.init = 16'h8000;
    LUT4 i7_3_lut (.A(\key_value[1] ), .B(\key_value[8] ), .C(\key_value[7] ), 
         .Z(n20_adj_821)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i7_3_lut.init = 16'h8080;
    LUT4 i9_4_lut (.A(\key_value[6] ), .B(\key_value[2] ), .C(\key_value[11] ), 
         .D(\key_value[3] ), .Z(n22_adj_823)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i9_4_lut.init = 16'h8000;
    LUT4 i3_2_lut (.A(\key_value[4] ), .B(\key_value[9] ), .Z(n16_adj_824)) /* synthesis lut_function=(A (B)) */ ;
    defparam i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_19 (.A(n3830), .B(n18679), .C(n436), .D(n18676), 
         .Z(\rom1_4__N_338[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_19.init = 16'hcfce;
    LUT4 i7545_4_lut (.A(n351), .B(n18763), .C(n18761), .D(n18771), 
         .Z(n414)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(65[4] 66[24])
    defparam i7545_4_lut.init = 16'hcfce;
    LUT4 i1_3_lut_4_lut_adj_20 (.A(n18684), .B(n18736), .C(n18735), .D(n18754), 
         .Z(n31)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A ((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(47[4] 48[25])
    defparam i1_3_lut_4_lut_adj_20.init = 16'h00f2;
    LUT4 i2_3_lut_4_lut_adj_21 (.A(n18707), .B(n18682), .C(n16888), .D(n18610), 
         .Z(clk_N_168_enable_514)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_21.init = 16'hfffe;
    CCU2D sub_6_add_2_9 (.A0(cycle[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cycle[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15309), 
          .COUT(n15310), .S0(CNT_17__N_703[7]), .S1(CNT_17__N_703[8]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_9.INIT0 = 16'h5555;
    defparam sub_6_add_2_9.INIT1 = 16'h5555;
    defparam sub_6_add_2_9.INJECT1_0 = "NO";
    defparam sub_6_add_2_9.INJECT1_1 = "NO";
    LUT4 i12286_3_lut (.A(n29), .B(n17345), .C(n30_adj_825), .Z(n15951)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(109[10:22])
    defparam i12286_3_lut.init = 16'h0404;
    LUT4 i11_4_lut_adj_22 (.A(CNT[13]), .B(CNT[7]), .C(CNT[8]), .D(CNT[12]), 
         .Z(n29)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(109[10:22])
    defparam i11_4_lut_adj_22.init = 16'hfffe;
    LUT4 i12285_4_lut (.A(n31_adj_826), .B(CNT[9]), .C(n28_adj_827), .D(CNT[2]), 
         .Z(n17345)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(109[10:22])
    defparam i12285_4_lut.init = 16'h0001;
    LUT4 i12_4_lut_adj_23 (.A(CNT[3]), .B(CNT[10]), .C(CNT[5]), .D(CNT[0]), 
         .Z(n30_adj_825)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(109[10:22])
    defparam i12_4_lut_adj_23.init = 16'hfffe;
    LUT4 i13_4_lut (.A(CNT[17]), .B(CNT[15]), .C(CNT[16]), .D(CNT[4]), 
         .Z(n31_adj_826)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(109[10:22])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(CNT[1]), .B(CNT[6]), .C(CNT[14]), .D(CNT[11]), 
         .Z(n28_adj_827)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(109[10:22])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i7439_2_lut (.A(n34), .B(CNT[17]), .Z(PWM_N_764)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i7439_2_lut.init = 16'h2222;
    LUT4 i7535_4_lut (.A(n247), .B(n18755), .C(n18708), .D(n18754), 
         .Z(n331)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(57[4] 58[25])
    defparam i7535_4_lut.init = 16'hcfce;
    LUT4 i9386_4_lut_then_4_lut (.A(\key_value[2] ), .B(\rom2[1] ), .C(n18721), 
         .D(\key_flag[2] ), .Z(n18849)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)+!B (C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(18[27:31])
    defparam i9386_4_lut_then_4_lut.init = 16'h7430;
    LUT4 i9386_4_lut_else_4_lut (.A(\key_flag[1] ), .B(\key_value[1] ), 
         .C(\rom2[1] ), .Z(n18848)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(18[27:31])
    defparam i9386_4_lut_else_4_lut.init = 16'h2020;
    LUT4 i1_2_lut_4_lut_adj_24 (.A(n16888), .B(n18623), .C(n18709), .D(n18648), 
         .Z(clk_N_168_enable_520)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_24.init = 16'hfffe;
    LUT4 i7474_2_lut_rep_552 (.A(\note[0] ), .B(\note[1] ), .Z(n18734)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(69[4] 88[14])
    defparam i7474_2_lut_rep_552.init = 16'hbbbb;
    LUT4 i12283_2_lut (.A(rst_n_c), .B(key_pa_c), .Z(pwm_out1_N_122)) /* synthesis lut_function=((B)+!A) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(25[10:16])
    defparam i12283_2_lut.init = 16'hdddd;
    CCU2D sub_6_add_2_7 (.A0(cycle[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cycle[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n15308), 
          .COUT(n15309), .S0(CNT_17__N_703[5]), .S1(CNT_17__N_703[6]));   // d:/fpga_project/lattice_diamond/piano/buzzer.v(27[19:28])
    defparam sub_6_add_2_7.INIT0 = 16'h5555;
    defparam sub_6_add_2_7.INIT1 = 16'h5555;
    defparam sub_6_add_2_7.INJECT1_0 = "NO";
    defparam sub_6_add_2_7.INJECT1_1 = "NO";
    LUT4 i4020_2_lut_3_lut_4_lut_4_lut (.A(yinjie[2]), .B(n19846), .C(n18785), 
         .D(n18784), .Z(n19839)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(29[9] 34[7])
    defparam i4020_2_lut_3_lut_4_lut_4_lut.init = 16'hd022;
    LUT4 i2_3_lut_4_lut_adj_25 (.A(n19846), .B(n18640), .C(n18610), .D(n18706), 
         .Z(clk_N_168_enable_522)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(55[4] 56[25])
    defparam i2_3_lut_4_lut_adj_25.init = 16'hfffe;
    LUT4 i1_2_lut_rep_435_3_lut_4_lut (.A(n18722), .B(n18682), .C(n19846), 
         .D(n18736), .Z(n18617)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(45[4] 46[25])
    defparam i1_2_lut_rep_435_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut_adj_26 (.A(n18684), .B(n18680), .C(n18706), .D(n18736), 
         .Z(n16876)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut_adj_26.init = 16'hfffe;
    LUT4 i5_4_lut (.A(n9), .B(n9654), .C(n8_adj_828), .D(n18722), .Z(clk_N_168_enable_508)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i5_4_lut.init = 16'hfffe;
    LUT4 i7541_4_lut (.A(n18725), .B(n18768), .C(n18755), .D(n10160), 
         .Z(n344)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B+!(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(59[4] 60[25])
    defparam i7541_4_lut.init = 16'hcfcd;
    LUT4 i11790_4_lut (.A(n18739), .B(n18749), .C(n18748), .D(n11), 
         .Z(n17081)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(111[11:24])
    defparam i11790_4_lut.init = 16'h5554;
    LUT4 i3_4_lut (.A(n18650), .B(n18754), .C(n18696), .D(n18606), .Z(clk_N_168_enable_509)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i3_4_lut_adj_27 (.A(n18612), .B(n18651), .C(n18763), .D(n18617), 
         .Z(clk_N_168_enable_510)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(55[4] 56[25])
    defparam i3_4_lut_adj_27.init = 16'hfffe;
    LUT4 i3_4_lut_adj_28 (.A(n18755), .B(n18640), .C(n18651), .D(n16920), 
         .Z(clk_N_168_enable_513)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(55[4] 56[25])
    defparam i3_4_lut_adj_28.init = 16'hfffe;
    LUT4 i3_4_lut_adj_29 (.A(n10337), .B(n18649), .C(n18685), .D(n16920), 
         .Z(clk_N_168_enable_515)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(45[4] 46[25])
    defparam i3_4_lut_adj_29.init = 16'hfffe;
    LUT4 i3_4_lut_adj_30 (.A(n18652), .B(n18755), .C(n10160), .D(n18619), 
         .Z(clk_N_168_enable_516)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(196[7] 205[5])
    defparam i3_4_lut_adj_30.init = 16'hfffe;
    LUT4 i4_4_lut (.A(n9654), .B(n16909), .C(n10160), .D(n6_adj_807), 
         .Z(clk_N_168_enable_517)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/buzzer.v(63[4] 64[24])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut_4_lut (.A(n18771), .B(n18709), .C(n18682), .D(n19846), 
         .Z(n8_adj_828)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module key_U17
//

module key_U17 (clk_N_168, \key_flag[4] , key_c_4, \key_value[4] , GND_net, 
            n18735, n6, n5, n891, n19846, n18754, n16888, n18747, 
            n5_adj_3, n11464, n18722, n18654, n18736, n312) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[4] ;
    input key_c_4;
    output \key_value[4] ;
    input GND_net;
    output n18735;
    input n6;
    input n5;
    output n891;
    input n19846;
    input n18754;
    output n16888;
    input n18747;
    input n5_adj_3;
    output n11464;
    input n18722;
    input n18654;
    input n18736;
    output n312;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18798, n10376, key_flag_N_639, key_reg, n15704;
    wire [31:0]n9;
    
    wire n15703, n15702, n15701, n15700, n15699, n15698, n15697, 
        n15696, n15695, n15694, n15693, n15692, n15691, n15690, 
        n15689, clk_N_168_enable_325, clk_N_168_enable_320;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n55, n60, n49, n50, n10219, n48, n39_adj_798, n58, 
        n52, n40_adj_799, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10376), .CK(clk_N_168), .CD(n18798), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[4] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_4), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_4), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[4] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15704), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15703), .COUT(n15704), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15702), .COUT(n15703), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15701), .COUT(n15702), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15700), .COUT(n15701), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15699), .COUT(n15700), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15698), .COUT(n15699), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15697), .COUT(n15698), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15696), .COUT(n15697), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15695), .COUT(n15696), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15694), .COUT(n15695), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15693), .COUT(n15694), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15692), .COUT(n15693), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15691), .COUT(n15692), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15690), .COUT(n15691), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15689), .COUT(n15690), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15689), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_320), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_325), .CD(n18798), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=82, LSE_RLINE=88 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10219)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_798), .B(n58), .C(n52), .D(n40_adj_799), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_798)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_799)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12281_2_lut (.A(delay_cnt[0]), .B(n10219), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12281_2_lut.init = 16'h2222;
    LUT4 key_reg_I_0_2_lut_rep_616 (.A(key_reg), .B(key_c_4), .Z(n18798)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_616.init = 16'h6666;
    LUT4 i7460_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7460_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7461_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7461_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7462_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7462_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7463_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7463_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7464_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7464_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7465_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7465_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_4), .C(n10219), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_320)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i7466_2_lut_3_lut (.A(key_reg), .B(key_c_4), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7466_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i5532_2_lut_rep_453 (.A(delay_cnt[0]), .B(n10219), .Z(clk_N_168_enable_325)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5532_2_lut_rep_453.init = 16'heeee;
    LUT4 i5533_2_lut_3_lut (.A(delay_cnt[0]), .B(n10219), .C(n9[0]), .Z(n10376)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5533_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_553 (.A(\key_flag[4] ), .B(\key_value[4] ), .Z(n18735)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_553.init = 16'h2222;
    LUT4 i289_3_lut_4_lut (.A(\key_flag[4] ), .B(\key_value[4] ), .C(n6), 
         .D(n5), .Z(n891)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i289_3_lut_4_lut.init = 16'h2220;
    LUT4 i1_2_lut_3_lut_4_lut_adj_16 (.A(\key_flag[4] ), .B(\key_value[4] ), 
         .C(n19846), .D(n18754), .Z(n16888)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_16.init = 16'hfff2;
    LUT4 i1_3_lut_4_lut (.A(\key_flag[4] ), .B(\key_value[4] ), .C(n18747), 
         .D(n5_adj_3), .Z(n11464)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2220;
    LUT4 i1_4_lut (.A(n18722), .B(n18654), .C(n18735), .D(n18736), .Z(n312)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i1_4_lut.init = 16'h3032;
    
endmodule
//
// Verilog Description of module key_U14
//

module key_U14 (clk_N_168, \key_flag[7] , key_c_7, \key_value[7] , GND_net, 
            n18756, n18770, n18758, n37, n34, \cycle_17__N_740[10] , 
            n19846, \cycle_17__N_663[10] , n18815, \key_flag[8] , \key_value[8] , 
            n18685, \key_flag[6] , \key_value[6] , n18708, n456, n3800, 
            n464, n3815) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[7] ;
    input key_c_7;
    output \key_value[7] ;
    input GND_net;
    output n18756;
    input n18770;
    input n18758;
    output n37;
    input n34;
    input \cycle_17__N_740[10] ;
    input n19846;
    output \cycle_17__N_663[10] ;
    output n18815;
    input \key_flag[8] ;
    input \key_value[8] ;
    output n18685;
    input \key_flag[6] ;
    input \key_value[6] ;
    output n18708;
    input n456;
    input n3800;
    input n464;
    output n3815;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18795, n10382, key_flag_N_639, key_reg, clk_N_168_enable_232;
    wire [31:0]n9;
    
    wire clk_N_168_enable_227;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15656, n15655, n15654, n15653, n15652, n15651, n15650, 
        n15649, n15648, n15647, n15646, n15645, n15644, n15643, 
        n15642, n15641, n10240, n55, n60, n49, n50, n48, n39_adj_796, 
        n58, n52, n40_adj_797, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10382), .CK(clk_N_168), .CD(n18795), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[7] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_7), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_7), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[7] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_227), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_232), .CD(n18795), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=107, LSE_RLINE=113 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15656), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15655), .COUT(n15656), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15654), .COUT(n15655), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15653), .COUT(n15654), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15652), .COUT(n15653), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15651), .COUT(n15652), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15650), .COUT(n15651), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15649), .COUT(n15650), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15648), .COUT(n15649), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15647), .COUT(n15648), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15646), .COUT(n15647), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15645), .COUT(n15646), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15644), .COUT(n15645), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15643), .COUT(n15644), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15642), .COUT(n15643), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15641), .COUT(n15642), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15641), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_574 (.A(\key_value[7] ), .B(\key_flag[7] ), .Z(n18756)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(12[17:25])
    defparam i1_2_lut_rep_574.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\key_value[7] ), .B(\key_flag[7] ), .C(n18770), 
         .D(n18758), .Z(n37)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(12[17:25])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hbbbf;
    LUT4 i5538_2_lut_rep_449 (.A(delay_cnt[0]), .B(n10240), .Z(clk_N_168_enable_232)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5538_2_lut_rep_449.init = 16'heeee;
    LUT4 i5539_2_lut_3_lut (.A(delay_cnt[0]), .B(n10240), .C(n9[0]), .Z(n10382)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5539_2_lut_3_lut.init = 16'he0e0;
    PFUMX i6554 (.BLUT(n34), .ALUT(\cycle_17__N_740[10] ), .C0(n19846), 
          .Z(\cycle_17__N_663[10] ));
    LUT4 key_reg_I_0_2_lut_rep_613 (.A(key_reg), .B(key_c_7), .Z(n18795)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_613.init = 16'h6666;
    LUT4 i7400_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7400_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7401_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7401_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7402_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7402_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7405_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7405_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7406_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7406_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7409_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7409_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7410_2_lut_3_lut (.A(key_reg), .B(key_c_7), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7410_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_15 (.A(key_reg), .B(key_c_7), .C(n10240), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_227)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut_adj_15.init = 16'hfff6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10240)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_796), .B(n58), .C(n52), .D(n40_adj_797), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_796)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_797)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12301_2_lut (.A(delay_cnt[0]), .B(n10240), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12301_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_633 (.A(\key_value[7] ), .B(\key_flag[7] ), .Z(n18815)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_633.init = 16'h4444;
    LUT4 i1_2_lut_rep_503_3_lut_4_lut (.A(\key_value[7] ), .B(\key_flag[7] ), 
         .C(\key_flag[8] ), .D(\key_value[8] ), .Z(n18685)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_503_3_lut_4_lut.init = 16'h44f4;
    LUT4 i1_2_lut_rep_526_3_lut_4_lut (.A(\key_value[7] ), .B(\key_flag[7] ), 
         .C(\key_flag[6] ), .D(\key_value[6] ), .Z(n18708)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_526_3_lut_4_lut.init = 16'h44f4;
    LUT4 i1_4_lut (.A(n456), .B(n37), .C(n3800), .D(n464), .Z(n3815)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(12[17:25])
    defparam i1_4_lut.init = 16'heeea;
    
endmodule
//
// Verilog Description of module key_U27
//

module key_U27 (GND_net, clk_N_168, \key_flag[9] , key_c_9, \key_value[9] , 
            n18768, \key_flag[8] , \key_value[8] , n9654, \rom2[0] , 
            n18771, n17235, n6, n5, n911) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk_N_168;
    output \key_flag[9] ;
    input key_c_9;
    output \key_value[9] ;
    output n18768;
    input \key_flag[8] ;
    input \key_value[8] ;
    output n9654;
    input \rom2[0] ;
    input n18771;
    output n17235;
    input n6;
    input n5;
    output n911;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15614;
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    wire [31:0]n9;
    
    wire n15615, n15613, n15612, n15611, n15610, n15609, n18793, 
        n10386, key_flag_N_639, key_reg, clk_N_168_enable_170, clk_N_168_enable_165;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n10246, n15624, n15623, n55, n60, n49, n50, n48, n39_adj_792, 
        n58, n52, n40_adj_793, n54, n44, n15622, n15621, n15620, 
        n15619, n15618, n15617, n15616;
    
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15614), .COUT(n15615), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15613), .COUT(n15614), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15612), .COUT(n15613), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15611), .COUT(n15612), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15610), .COUT(n15611), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15609), .COUT(n15610), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15609), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    FD1S3IX delay_cnt_i0 (.D(n10386), .CK(clk_N_168), .CD(n18793), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[9] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_9), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_9), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[9] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_165), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_170), .CD(n18793), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=124, LSE_RLINE=130 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i5542_2_lut_rep_447 (.A(delay_cnt[0]), .B(n10246), .Z(clk_N_168_enable_170)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5542_2_lut_rep_447.init = 16'heeee;
    LUT4 i5543_2_lut_3_lut (.A(delay_cnt[0]), .B(n10246), .C(n9[0]), .Z(n10386)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5543_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_586 (.A(\key_flag[9] ), .B(\key_value[9] ), .Z(n18768)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_586.init = 16'h2222;
    LUT4 i4_2_lut_3_lut_4_lut (.A(\key_flag[9] ), .B(\key_value[9] ), .C(\key_flag[8] ), 
         .D(\key_value[8] ), .Z(n9654)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i4_2_lut_3_lut_4_lut.init = 16'h22f2;
    LUT4 i11944_3_lut_4_lut (.A(\key_flag[9] ), .B(\key_value[9] ), .C(\rom2[0] ), 
         .D(n18771), .Z(n17235)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i11944_3_lut_4_lut.init = 16'hf202;
    LUT4 i309_3_lut_4_lut (.A(\key_flag[9] ), .B(\key_value[9] ), .C(n6), 
         .D(n5), .Z(n911)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i309_3_lut_4_lut.init = 16'h2220;
    LUT4 key_reg_I_0_2_lut_rep_611 (.A(key_reg), .B(key_c_9), .Z(n18793)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_611.init = 16'h6666;
    LUT4 i7374_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7374_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7375_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7375_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7376_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7376_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7377_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7377_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7378_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7378_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7379_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7379_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7380_2_lut_3_lut (.A(key_reg), .B(key_c_9), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7380_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_9), .C(n10246), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_165)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15624), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15623), .COUT(n15624), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10246)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_792), .B(n58), .C(n52), .D(n40_adj_793), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_792)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_793)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12305_2_lut (.A(delay_cnt[0]), .B(n10246), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12305_2_lut.init = 16'h2222;
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15622), .COUT(n15623), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15621), .COUT(n15622), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15620), .COUT(n15621), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15619), .COUT(n15620), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15618), .COUT(n15619), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15617), .COUT(n15618), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15616), .COUT(n15617), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15615), .COUT(n15616), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module key_U26
//

module key_U26 (clk_N_168, \key_flag[10] , key_c_10, \key_value[10] , 
            GND_net, n18771, n18761, n344, n18763, n407, n9654, 
            n312, n18709, n417, n18768, n321, n405, \key_flag[11] , 
            \key_value[11] , n16909, n6, n18813, n18719, \key_value[9] , 
            \key_flag[9] , n18667) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[10] ;
    input key_c_10;
    output \key_value[10] ;
    input GND_net;
    output n18771;
    input n18761;
    input n344;
    input n18763;
    output n407;
    input n9654;
    input n312;
    input n18709;
    output n417;
    input n18768;
    input n321;
    output n405;
    input \key_flag[11] ;
    input \key_value[11] ;
    output n16909;
    input n6;
    input n18813;
    output n18719;
    input \key_value[9] ;
    input \key_flag[9] ;
    output n18667;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18792, n10388, key_flag_N_639, key_reg, n15608;
    wire [31:0]n9;
    
    wire n15607, n15606, n15605, n15604, n15603, n15602, n15601, 
        n15600, n15599, n15598, n15597, n15596, n15595, n15594, 
        n15593, clk_N_168_enable_139, clk_N_168_enable_134;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n10249, n55, n60, n49, n50, n48, n39_adj_790, n58, 
        n52, n40_adj_791, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10388), .CK(clk_N_168), .CD(n18792), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[10] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_10), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_10), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[10] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15608), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15607), .COUT(n15608), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15606), .COUT(n15607), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15605), .COUT(n15606), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15604), .COUT(n15605), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15603), .COUT(n15604), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15602), .COUT(n15603), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15601), .COUT(n15602), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15600), .COUT(n15601), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15599), .COUT(n15600), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15598), .COUT(n15599), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15597), .COUT(n15598), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15596), .COUT(n15597), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15595), .COUT(n15596), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15594), .COUT(n15595), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15593), .COUT(n15594), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15593), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_134), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_139), .CD(n18792), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=132, LSE_RLINE=138 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i7548_4_lut_4_lut_4_lut (.A(n18771), .B(n18761), .C(n344), .D(n18763), 
         .Z(n407)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i7548_4_lut_4_lut_4_lut.init = 16'h00dc;
    LUT4 i8055_4_lut_4_lut (.A(n18771), .B(n9654), .C(n312), .D(n18709), 
         .Z(n417)) /* synthesis lut_function=(A (D)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i8055_4_lut_4_lut.init = 16'hff54;
    LUT4 i8052_4_lut_4_lut (.A(n18771), .B(n18768), .C(n321), .D(n18709), 
         .Z(n405)) /* synthesis lut_function=(A (D)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i8052_4_lut_4_lut.init = 16'hff54;
    LUT4 i5544_2_lut_rep_446 (.A(delay_cnt[0]), .B(n10249), .Z(clk_N_168_enable_139)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5544_2_lut_rep_446.init = 16'heeee;
    LUT4 i5545_2_lut_3_lut (.A(delay_cnt[0]), .B(n10249), .C(n9[0]), .Z(n10388)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5545_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_589 (.A(\key_value[10] ), .B(\key_flag[10] ), .Z(n18771)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_589.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\key_value[10] ), .B(\key_flag[10] ), 
         .C(\key_flag[11] ), .D(\key_value[11] ), .Z(n16909)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h44f4;
    LUT4 i313_3_lut_rep_537_4_lut (.A(\key_value[10] ), .B(\key_flag[10] ), 
         .C(n6), .D(n18813), .Z(n18719)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i313_3_lut_rep_537_4_lut.init = 16'h4044;
    LUT4 i12314_2_lut_rep_485_2_lut_3_lut_4_lut (.A(\key_value[10] ), .B(\key_flag[10] ), 
         .C(\key_value[9] ), .D(\key_flag[9] ), .Z(n18667)) /* synthesis lut_function=(A (C+!(D))+!A !(B+!(C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i12314_2_lut_rep_485_2_lut_3_lut_4_lut.init = 16'hb0bb;
    LUT4 key_reg_I_0_2_lut_rep_610 (.A(key_reg), .B(key_c_10), .Z(n18792)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_610.init = 16'h6666;
    LUT4 i7366_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7366_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7367_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7367_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7368_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7368_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7369_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7369_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7370_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7370_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7371_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7371_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7372_2_lut_3_lut (.A(key_reg), .B(key_c_10), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7372_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_14 (.A(key_reg), .B(key_c_10), .C(n10249), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_134)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut_adj_14.init = 16'hfff6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10249)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_790), .B(n58), .C(n52), .D(n40_adj_791), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_790)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_791)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12307_2_lut (.A(delay_cnt[0]), .B(n10249), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12307_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module key_U25
//

module key_U25 (clk_N_168, \key_flag[11] , key_c_11, \key_value[11] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[11] ;
    input key_c_11;
    output \key_value[11] ;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18791, n10390, key_flag_N_639, key_reg, clk_N_168_enable_108;
    wire [31:0]n9;
    
    wire n15592, n15591, n15590, n15589, n15588, n15587, n15586, 
        n15585, clk_N_168_enable_103;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15584, n15583, n15582, n15581, n15580, n15579, n15578, 
        n15577, n10252, n55, n60, n49, n50, n48, n39_adj_788, 
        n58, n52, n40_adj_789, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10390), .CK(clk_N_168), .CD(n18791), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[11] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_11), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_11), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[11] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15592), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15591), .COUT(n15592), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15590), .COUT(n15591), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15589), .COUT(n15590), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15588), .COUT(n15589), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15587), .COUT(n15588), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15586), .COUT(n15587), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15585), .COUT(n15586), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15584), .COUT(n15585), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15583), .COUT(n15584), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_103), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_108), .CD(n18791), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=140, LSE_RLINE=146 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15582), .COUT(n15583), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15581), .COUT(n15582), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15580), .COUT(n15581), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15579), .COUT(n15580), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15578), .COUT(n15579), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15577), .COUT(n15578), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15577), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i5546_2_lut_rep_445 (.A(delay_cnt[0]), .B(n10252), .Z(clk_N_168_enable_108)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5546_2_lut_rep_445.init = 16'heeee;
    LUT4 i5547_2_lut_3_lut (.A(delay_cnt[0]), .B(n10252), .C(n9[0]), .Z(n10390)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5547_2_lut_3_lut.init = 16'he0e0;
    LUT4 key_reg_I_0_2_lut_rep_609 (.A(key_reg), .B(key_c_11), .Z(n18791)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_609.init = 16'h6666;
    LUT4 i7359_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7359_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7360_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7360_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7361_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7361_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7362_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7362_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7363_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7363_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7364_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7364_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7365_2_lut_3_lut (.A(key_reg), .B(key_c_11), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7365_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_11), .C(n10252), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_103)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10252)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_788), .B(n58), .C(n52), .D(n40_adj_789), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_788)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_789)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12316_2_lut (.A(delay_cnt[0]), .B(n10252), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12316_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module key_U20
//

module key_U20 (clk_N_168, \key_flag[1] , key_c_1, \key_value[1] , GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[1] ;
    input key_c_1;
    output \key_value[1] ;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18801, n10370, key_flag_N_639, key_reg, n15363;
    wire [31:0]n9;
    
    wire n15362, n15361, n15360, n15359, n15358, n15357, n15356, 
        n15355, n15354, n15353, n15352, n15351, n15350, n15349, 
        n15348, clk_N_168_enable_419, clk_N_168_enable_414;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n55, n60, n49, n50, n10228, n48, n39_adj_786, n58, 
        n52, n40_adj_787, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10370), .CK(clk_N_168), .CD(n18801), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[1] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_1), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_1), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[1] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15363), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15362), .COUT(n15363), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15361), .COUT(n15362), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15360), .COUT(n15361), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15359), .COUT(n15360), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15358), .COUT(n15359), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15357), .COUT(n15358), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15356), .COUT(n15357), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15355), .COUT(n15356), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15354), .COUT(n15355), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15353), .COUT(n15354), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15352), .COUT(n15353), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15351), .COUT(n15352), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15350), .COUT(n15351), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15349), .COUT(n15350), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15348), .COUT(n15349), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15348), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_414), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_419), .CD(n18801), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=57, LSE_RLINE=63 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10228)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_786), .B(n58), .C(n52), .D(n40_adj_787), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_786)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_787)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12293_2_lut (.A(delay_cnt[0]), .B(n10228), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12293_2_lut.init = 16'h2222;
    LUT4 key_reg_I_0_2_lut_rep_619 (.A(key_reg), .B(key_c_1), .Z(n18801)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_619.init = 16'h6666;
    LUT4 i7495_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7495_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7496_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7496_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7497_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7497_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7498_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7498_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7499_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7499_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7500_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7500_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_1), .C(n10228), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_414)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i7501_2_lut_3_lut (.A(key_reg), .B(key_c_1), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7501_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i5526_2_lut_rep_456 (.A(delay_cnt[0]), .B(n10228), .Z(clk_N_168_enable_419)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5526_2_lut_rep_456.init = 16'heeee;
    LUT4 i5527_2_lut_3_lut (.A(delay_cnt[0]), .B(n10228), .C(n9[0]), .Z(n10370)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5527_2_lut_3_lut.init = 16'he0e0;
    
endmodule
//
// Verilog Description of module key_U24
//

module key_U24 (clk_N_168, \key_flag[12] , key_c_12, \key_value[12] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[12] ;
    input key_c_12;
    output \key_value[12] ;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18790, n10392, key_flag_N_639, key_reg, clk_N_168_enable_77;
    wire [31:0]n9;
    
    wire clk_N_168_enable_72;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15576, n15575, n15574, n15573, n15572, n15571, n15570, 
        n15569, n15568, n15567, n15566, n15565, n15564, n15563, 
        n15562, n15561, n10255, n55, n60, n49, n50, n48, n39_adj_784, 
        n58, n52, n40_adj_785, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10392), .CK(clk_N_168), .CD(n18790), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[12] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_12), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_12), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[12] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_72), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_77), .CD(n18790), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=148, LSE_RLINE=154 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15576), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15575), .COUT(n15576), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15574), .COUT(n15575), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15573), .COUT(n15574), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15572), .COUT(n15573), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15571), .COUT(n15572), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15570), .COUT(n15571), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15569), .COUT(n15570), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15568), .COUT(n15569), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15567), .COUT(n15568), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15566), .COUT(n15567), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15565), .COUT(n15566), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15564), .COUT(n15565), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15563), .COUT(n15564), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15562), .COUT(n15563), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15561), .COUT(n15562), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15561), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i5548_2_lut_rep_444 (.A(delay_cnt[0]), .B(n10255), .Z(clk_N_168_enable_77)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5548_2_lut_rep_444.init = 16'heeee;
    LUT4 i5549_2_lut_3_lut (.A(delay_cnt[0]), .B(n10255), .C(n9[0]), .Z(n10392)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5549_2_lut_3_lut.init = 16'he0e0;
    LUT4 key_reg_I_0_2_lut_rep_608 (.A(key_reg), .B(key_c_12), .Z(n18790)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_608.init = 16'h6666;
    LUT4 i7354_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7354_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7353_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7353_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7352_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7352_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7351_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7351_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7350_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7350_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7355_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7355_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7358_2_lut_3_lut (.A(key_reg), .B(key_c_12), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7358_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_12), .C(n10255), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_72)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10255)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_784), .B(n58), .C(n52), .D(n40_adj_785), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_784)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_785)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12318_2_lut (.A(delay_cnt[0]), .B(n10255), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12318_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module key_U13
//

module key_U13 (clk_N_168, \key_flag[8] , key_c_8, \key_value[8] , GND_net, 
            n18755, \rom2[0] , n18815, n17234, n18770, n5, n464, 
            n6, n5_adj_2, n907, n18768, n16917) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[8] ;
    input key_c_8;
    output \key_value[8] ;
    input GND_net;
    output n18755;
    input \rom2[0] ;
    input n18815;
    output n17234;
    input n18770;
    input n5;
    output n464;
    input n6;
    input n5_adj_2;
    output n907;
    input n18768;
    output n16917;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18794, n10384, key_flag_N_639, key_reg, clk_N_168_enable_201;
    wire [31:0]n9;
    
    wire clk_N_168_enable_196;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15640, n15639, n15638, n15637, n15636, n15635, n15634, 
        n15633, n15632, n10243, n15631, n15630, n15629, n15628, 
        n15627, n15626, n15625, n55, n60, n49, n50, n48, n39_adj_782, 
        n58, n52, n40_adj_783, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10384), .CK(clk_N_168), .CD(n18794), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[8] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_8), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_8), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[8] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_196), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_201), .CD(n18794), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=116, LSE_RLINE=122 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15640), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15639), .COUT(n15640), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15638), .COUT(n15639), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15637), .COUT(n15638), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15636), .COUT(n15637), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15635), .COUT(n15636), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15634), .COUT(n15635), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15633), .COUT(n15634), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15632), .COUT(n15633), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_573 (.A(\key_value[8] ), .B(\key_flag[8] ), .Z(n18755)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_573.init = 16'h4444;
    LUT4 i11943_3_lut_4_lut (.A(\key_value[8] ), .B(\key_flag[8] ), .C(\rom2[0] ), 
         .D(n18815), .Z(n17234)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i11943_3_lut_4_lut.init = 16'h4f40;
    LUT4 i117_3_lut_4_lut (.A(\key_value[8] ), .B(\key_flag[8] ), .C(n18770), 
         .D(n5), .Z(n464)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i117_3_lut_4_lut.init = 16'h4440;
    LUT4 i305_3_lut_4_lut (.A(\key_value[8] ), .B(\key_flag[8] ), .C(n6), 
         .D(n5_adj_2), .Z(n907)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i305_3_lut_4_lut.init = 16'h4440;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\key_value[8] ), .B(\key_flag[8] ), .C(n18768), 
         .D(n18815), .Z(n16917)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i5540_2_lut_rep_448 (.A(delay_cnt[0]), .B(n10243), .Z(clk_N_168_enable_201)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5540_2_lut_rep_448.init = 16'heeee;
    LUT4 i5541_2_lut_3_lut (.A(delay_cnt[0]), .B(n10243), .C(n9[0]), .Z(n10384)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5541_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15631), .COUT(n15632), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15630), .COUT(n15631), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15629), .COUT(n15630), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15628), .COUT(n15629), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15627), .COUT(n15628), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15626), .COUT(n15627), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    LUT4 key_reg_I_0_2_lut_rep_612 (.A(key_reg), .B(key_c_8), .Z(n18794)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_612.init = 16'h6666;
    LUT4 i7387_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7387_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7390_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7390_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7391_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7391_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7385_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7385_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7386_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7386_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7392_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7392_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7393_2_lut_3_lut (.A(key_reg), .B(key_c_8), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7393_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut_adj_13 (.A(key_reg), .B(key_c_8), .C(n10243), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_196)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut_adj_13.init = 16'hfff6;
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15625), .COUT(n15626), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15625), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10243)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_782), .B(n58), .C(n52), .D(n40_adj_783), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_782)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_783)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12303_2_lut (.A(delay_cnt[0]), .B(n10243), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12303_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module key_U21
//

module key_U21 (GND_net, \key_value[0] , clk_N_168, key_c_0, \key_flag[0] , 
            n5, n18721, n18724, n9292, n18644, n6, n5_adj_1, n18713, 
            n19846, n18680, n18679, n18722, n18725, n18649, n18652) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \key_value[0] ;
    input clk_N_168;
    input key_c_0;
    output \key_flag[0] ;
    input n5;
    output n18721;
    input n18724;
    input n9292;
    output n18644;
    input n6;
    input n5_adj_1;
    output n18713;
    input n19846;
    output n18680;
    output n18679;
    input n18722;
    input n18725;
    output n18649;
    output n18652;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    wire n15371;
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    wire [31:0]n9;
    
    wire n15372, key_flag_N_639, n18802, n10368, key_reg, n15370, 
        n15369, n15368, n15367, n15366, n15365, n15364, clk_N_168_enable_450, 
        clk_N_168_enable_445;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n10222, n55, n60, n49, n50, n48, n39_adj_778, n58, 
        n52, n40_adj_779, n54, n44, n15379, n15378, n15377, n15376, 
        n15375, n15374, n15373;
    
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15371), .COUT(n15372), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    FD1P3AY key_value_28 (.D(key_c_0), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[0] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1S3IX delay_cnt_i0 (.D(n10368), .CK(clk_N_168), .CD(n18802), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[0] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_0), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15370), .COUT(n15371), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15369), .COUT(n15370), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15368), .COUT(n15369), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15367), .COUT(n15368), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15366), .COUT(n15367), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15365), .COUT(n15366), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15364), .COUT(n15365), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15364), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_462_4_lut (.A(n5), .B(n18721), .C(n18724), .D(n9292), 
         .Z(n18644)) /* synthesis lut_function=(A (B+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_462_4_lut.init = 16'hffc8;
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_445), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_450), .CD(n18802), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=48, LSE_RLINE=54 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i12265_2_lut (.A(delay_cnt[0]), .B(n10222), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12265_2_lut.init = 16'h2222;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10222)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_778), .B(n58), .C(n52), .D(n40_adj_779), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_778)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_779)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13_2_lut.init = 16'heeee;
    LUT4 key_reg_I_0_2_lut_rep_620 (.A(key_reg), .B(key_c_0), .Z(n18802)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_620.init = 16'h6666;
    LUT4 i7503_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7503_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7504_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7504_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7505_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7505_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7506_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7506_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7507_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7507_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7508_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7508_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_0), .C(n10222), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_445)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i7509_2_lut_3_lut (.A(key_reg), .B(key_c_0), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7509_2_lut_3_lut.init = 16'hf6f6;
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15379), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15378), .COUT(n15379), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15377), .COUT(n15378), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    LUT4 i5524_2_lut_rep_457 (.A(delay_cnt[0]), .B(n10222), .Z(clk_N_168_enable_450)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5524_2_lut_rep_457.init = 16'heeee;
    LUT4 i5525_2_lut_3_lut (.A(delay_cnt[0]), .B(n10222), .C(n9[0]), .Z(n10368)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5525_2_lut_3_lut.init = 16'he0e0;
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15376), .COUT(n15377), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15375), .COUT(n15376), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_539 (.A(\key_value[0] ), .B(\key_flag[0] ), .Z(n18721)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_539.init = 16'h4444;
    LUT4 i273_3_lut_rep_531_4_lut (.A(\key_value[0] ), .B(\key_flag[0] ), 
         .C(n6), .D(n5_adj_1), .Z(n18713)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i273_3_lut_rep_531_4_lut.init = 16'h4440;
    LUT4 i1_2_lut_rep_498_3_lut (.A(\key_value[0] ), .B(\key_flag[0] ), 
         .C(n19846), .Z(n18680)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_498_3_lut.init = 16'hf4f4;
    LUT4 i1_3_lut_rep_497_4_lut (.A(\key_value[0] ), .B(\key_flag[0] ), 
         .C(n18724), .D(n5), .Z(n18679)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_3_lut_rep_497_4_lut.init = 16'h4440;
    LUT4 i2_2_lut_rep_467_3_lut_4_lut (.A(\key_value[0] ), .B(\key_flag[0] ), 
         .C(n18722), .D(n18725), .Z(n18649)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i2_2_lut_rep_467_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_470_3_lut_4_lut (.A(\key_value[0] ), .B(\key_flag[0] ), 
         .C(n19846), .D(n18725), .Z(n18652)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_470_3_lut_4_lut.init = 16'hfff4;
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15374), .COUT(n15375), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15373), .COUT(n15374), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15372), .COUT(n15373), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module key_U15
//

module key_U15 (clk_N_168, \key_flag[6] , key_c_6, \key_value[6] , GND_net, 
            n18720, n18754, n18815, n18654, n18735, n18655, n6, 
            n18813, n18677, n18747, n12156, n456, \rom2[1] , n18597, 
            n18755, n18668) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[6] ;
    input key_c_6;
    output \key_value[6] ;
    input GND_net;
    output n18720;
    input n18754;
    input n18815;
    output n18654;
    input n18735;
    output n18655;
    input n6;
    input n18813;
    output n18677;
    input n18747;
    input n12156;
    output n456;
    input \rom2[1] ;
    output n18597;
    input n18755;
    output n18668;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18796, n10380, key_flag_N_639, key_reg, clk_N_168_enable_263;
    wire [31:0]n9;
    
    wire clk_N_168_enable_258;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15672, n15671, n15670, n15669, n15668, n15667, n15666, 
        n15665, n15664, n15663, n15662, n15661, n15660, n15659, 
        n15658, n15657, n10237, n55, n60, n49, n50, n48, n39_adj_776, 
        n58, n52, n40_adj_777, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10380), .CK(clk_N_168), .CD(n18796), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[6] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_6), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_6), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[6] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_258), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_263), .CD(n18796), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=98, LSE_RLINE=104 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15672), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15671), .COUT(n15672), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15670), .COUT(n15671), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15669), .COUT(n15670), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15668), .COUT(n15669), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15667), .COUT(n15668), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15666), .COUT(n15667), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15665), .COUT(n15666), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15664), .COUT(n15665), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15663), .COUT(n15664), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15662), .COUT(n15663), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15661), .COUT(n15662), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15660), .COUT(n15661), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15659), .COUT(n15660), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15658), .COUT(n15659), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15657), .COUT(n15658), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15657), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i5536_2_lut_rep_450 (.A(delay_cnt[0]), .B(n10237), .Z(clk_N_168_enable_263)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5536_2_lut_rep_450.init = 16'heeee;
    LUT4 i5537_2_lut_3_lut (.A(delay_cnt[0]), .B(n10237), .C(n9[0]), .Z(n10380)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5537_2_lut_3_lut.init = 16'he0e0;
    LUT4 key_reg_I_0_2_lut_rep_614 (.A(key_reg), .B(key_c_6), .Z(n18796)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_614.init = 16'h6666;
    LUT4 i7432_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7432_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7428_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7428_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7429_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7429_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7430_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7430_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7431_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7431_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7433_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7433_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7434_2_lut_3_lut (.A(key_reg), .B(key_c_6), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7434_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_6), .C(n10237), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_258)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10237)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_776), .B(n58), .C(n52), .D(n40_adj_777), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_776)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_777)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12299_2_lut (.A(delay_cnt[0]), .B(n10237), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12299_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_rep_538 (.A(\key_value[6] ), .B(\key_flag[6] ), .Z(n18720)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_538.init = 16'h4444;
    LUT4 i1_2_lut_rep_472_3_lut_4_lut (.A(\key_value[6] ), .B(\key_flag[6] ), 
         .C(n18754), .D(n18815), .Z(n18654)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_472_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_473_3_lut_4_lut (.A(\key_value[6] ), .B(\key_flag[6] ), 
         .C(n18735), .D(n18754), .Z(n18655)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_473_3_lut_4_lut.init = 16'hfff4;
    LUT4 i297_3_lut_rep_495_4_lut (.A(\key_value[6] ), .B(\key_flag[6] ), 
         .C(n6), .D(n18813), .Z(n18677)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i297_3_lut_rep_495_4_lut.init = 16'h4044;
    LUT4 i109_3_lut_4_lut (.A(\key_value[6] ), .B(\key_flag[6] ), .C(n18747), 
         .D(n12156), .Z(n456)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i109_3_lut_4_lut.init = 16'h4044;
    LUT4 n446_bdd_3_lut_12599_4_lut (.A(\key_value[6] ), .B(\key_flag[6] ), 
         .C(\rom2[1] ), .D(n18735), .Z(n18597)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam n446_bdd_3_lut_12599_4_lut.init = 16'h4f40;
    LUT4 i1_2_lut_rep_486_3_lut_4_lut (.A(\key_value[6] ), .B(\key_flag[6] ), 
         .C(n18755), .D(n18815), .Z(n18668)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_486_3_lut_4_lut.init = 16'hfff4;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module key_U16
//

module key_U16 (clk_N_168, \key_flag[5] , key_c_5, \key_value[5] , GND_net, 
            n18754, \key_value[4] , \key_flag[4] , n18706, n6, n5, 
            n895) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[5] ;
    input key_c_5;
    output \key_value[5] ;
    input GND_net;
    output n18754;
    input \key_value[4] ;
    input \key_flag[4] ;
    output n18706;
    input n6;
    input n5;
    output n895;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18797, n10378, key_flag_N_639, key_reg, n15688;
    wire [31:0]n9;
    
    wire n15687, n15686, n15685, n15684, n15683, n15682, n15681, 
        n15680, n15679, n15678, n15677, n15676, n15675, n15674, 
        n15673, clk_N_168_enable_294, clk_N_168_enable_289;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n10231, n55, n60, n49, n50, n48, n39_adj_774, n58, 
        n52, n40_adj_775, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10378), .CK(clk_N_168), .CD(n18797), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[5] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_5), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_5), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[5] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15688), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15687), .COUT(n15688), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15686), .COUT(n15687), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15685), .COUT(n15686), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15684), .COUT(n15685), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15683), .COUT(n15684), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15682), .COUT(n15683), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15681), .COUT(n15682), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15680), .COUT(n15681), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15679), .COUT(n15680), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15678), .COUT(n15679), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15677), .COUT(n15678), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15676), .COUT(n15677), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15675), .COUT(n15676), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15674), .COUT(n15675), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15673), .COUT(n15674), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15673), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_289), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_294), .CD(n18797), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=90, LSE_RLINE=96 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_572 (.A(\key_flag[5] ), .B(\key_value[5] ), .Z(n18754)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_572.init = 16'h2222;
    LUT4 i1_2_lut_rep_524_3_lut_4_lut (.A(\key_flag[5] ), .B(\key_value[5] ), 
         .C(\key_value[4] ), .D(\key_flag[4] ), .Z(n18706)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_524_3_lut_4_lut.init = 16'h2f22;
    LUT4 i293_3_lut_4_lut (.A(\key_flag[5] ), .B(\key_value[5] ), .C(n6), 
         .D(n5), .Z(n895)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i293_3_lut_4_lut.init = 16'h2220;
    LUT4 i5534_2_lut_rep_451 (.A(delay_cnt[0]), .B(n10231), .Z(clk_N_168_enable_294)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5534_2_lut_rep_451.init = 16'heeee;
    LUT4 i5535_2_lut_3_lut (.A(delay_cnt[0]), .B(n10231), .C(n9[0]), .Z(n10378)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5535_2_lut_3_lut.init = 16'he0e0;
    LUT4 key_reg_I_0_2_lut_rep_615 (.A(key_reg), .B(key_c_5), .Z(n18797)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_615.init = 16'h6666;
    LUT4 i7442_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7442_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7443_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7443_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7444_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7444_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7447_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7447_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7448_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7448_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7451_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7451_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_5), .C(n10231), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_289)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i7452_2_lut_3_lut (.A(key_reg), .B(key_c_5), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7452_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10231)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_774), .B(n58), .C(n52), .D(n40_adj_775), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_774)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_775)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12297_2_lut (.A(delay_cnt[0]), .B(n10231), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12297_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module key_U19
//

module key_U19 (clk_N_168, \key_flag[2] , key_c_2, \key_value[2] , GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[2] ;
    input key_c_2;
    output \key_value[2] ;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18800, n10372, key_flag_N_639, key_reg;
    wire [31:0]n9;
    
    wire n15332, n15333, n15347, n15346, n15345, n15344, n15343, 
        n15342, n15341, n15340, n15339, n15338, n15337, n15336, 
        n15335, n15334, clk_N_168_enable_387, clk_N_168_enable_382;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n55, n60, n49, n50, n10234, n48, n39_adj_772, n58, 
        n52, n40_adj_773, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10372), .CK(clk_N_168), .CD(n18800), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[2] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_2), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_2), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[2] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15332), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15332), .COUT(n15333), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15347), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15346), .COUT(n15347), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15345), .COUT(n15346), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15344), .COUT(n15345), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15343), .COUT(n15344), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15342), .COUT(n15343), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15341), .COUT(n15342), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15340), .COUT(n15341), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15339), .COUT(n15340), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15338), .COUT(n15339), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15337), .COUT(n15338), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15336), .COUT(n15337), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15335), .COUT(n15336), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15334), .COUT(n15335), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15333), .COUT(n15334), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_382), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_387), .CD(n18800), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=66, LSE_RLINE=72 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10234)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_772), .B(n58), .C(n52), .D(n40_adj_773), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_772)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_773)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12295_2_lut (.A(delay_cnt[0]), .B(n10234), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12295_2_lut.init = 16'h2222;
    LUT4 key_reg_I_0_2_lut_rep_618 (.A(key_reg), .B(key_c_2), .Z(n18800)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_618.init = 16'h6666;
    LUT4 i7487_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7487_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7488_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7488_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7489_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7489_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7490_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7490_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7491_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7491_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7492_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7492_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7494_2_lut_3_lut (.A(key_reg), .B(key_c_2), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7494_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_2), .C(n10234), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_382)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i5528_2_lut_rep_455 (.A(delay_cnt[0]), .B(n10234), .Z(clk_N_168_enable_387)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5528_2_lut_rep_455.init = 16'heeee;
    LUT4 i5529_2_lut_3_lut (.A(delay_cnt[0]), .B(n10234), .C(n9[0]), .Z(n10372)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5529_2_lut_3_lut.init = 16'he0e0;
    
endmodule
//
// Verilog Description of module key_U22
//

module key_U22 (clk_N_168, \key_flag[14] , key_c_14, \key_value[14] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[14] ;
    input key_c_14;
    output \key_value[14] ;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire clk_N_168_enable_462;
    wire [31:0]delay_cnt_31__N_570;
    
    wire clk_N_168_enable_531, n18728;
    wire [31:0]n9;
    
    wire n10396, key_flag_N_639, key_reg, n15544, n15543, n15542, 
        n15541, n15540, n15539, n15538, n15537, n15536, n15535, 
        n15534, n15533, n15532, n15531, n15530, n15529, n10261, 
        n55, n60, n49, n50, n48, n39_adj_770, n58, n52, n40_adj_771, 
        n54, n44;
    
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    FD1S3IX delay_cnt_i0 (.D(n10396), .CK(clk_N_168), .CD(n18728), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[14] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_14), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_14), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[14] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15544), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15543), .COUT(n15544), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15542), .COUT(n15543), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15541), .COUT(n15542), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15540), .COUT(n15541), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15539), .COUT(n15540), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15538), .COUT(n15539), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15537), .COUT(n15538), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15536), .COUT(n15537), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15535), .COUT(n15536), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15534), .COUT(n15535), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15533), .COUT(n15534), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15532), .COUT(n15533), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15531), .COUT(n15532), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15530), .COUT(n15531), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15529), .COUT(n15530), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15529), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i5553_2_lut_3_lut (.A(delay_cnt[0]), .B(n10261), .C(n9[0]), .Z(n10396)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5553_2_lut_3_lut.init = 16'he0e0;
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_462), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    LUT4 i12322_2_lut (.A(delay_cnt[0]), .B(n10261), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12322_2_lut.init = 16'h2222;
    LUT4 key_reg_I_0_2_lut_rep_546 (.A(key_reg), .B(key_c_14), .Z(n18728)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_546.init = 16'h6666;
    LUT4 i7298_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7298_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7301_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7301_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7300_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7300_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7307_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7307_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7306_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7306_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7299_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7299_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7297_2_lut_3_lut (.A(key_reg), .B(key_c_14), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7297_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_14), .C(n10261), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_462)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_531), .CD(n18728), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=164, LSE_RLINE=170 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10261)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_770), .B(n58), .C(n52), .D(n40_adj_771), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i5552_2_lut_rep_436 (.A(delay_cnt[0]), .B(n10261), .Z(clk_N_168_enable_531)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5552_2_lut_rep_436.init = 16'heeee;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_770)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_771)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module key_U18
//

module key_U18 (clk_N_168, \key_flag[3] , key_c_3, \key_value[3] , GND_net, 
            n18736, n6, n18814, n887, \rom2[1] , n18754, n18598, 
            \key_flag[2] , \key_value[2] , n18707, n18747, n18758, 
            n444, \key_value[4] , \key_flag[4] , n18696) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[3] ;
    input key_c_3;
    output \key_value[3] ;
    input GND_net;
    output n18736;
    input n6;
    input n18814;
    output n887;
    input \rom2[1] ;
    input n18754;
    output n18598;
    input \key_flag[2] ;
    input \key_value[2] ;
    output n18707;
    input n18747;
    input n18758;
    output n444;
    input \key_value[4] ;
    input \key_flag[4] ;
    output n18696;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18799, n10374, key_flag_N_639, key_reg, n15331;
    wire [31:0]n9;
    
    wire n15330, n15329, n15328, n15327, n15326, n15325, n15324, 
        n15323, n15322, n15321, n15320, n15319, n15318, clk_N_168_enable_356, 
        clk_N_168_enable_351;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15317, n55, n60, n49, n50, n10225, n48, n39_adj_768, 
        n58, n52, n40_adj_769, n54, n44, n15316;
    
    FD1S3IX delay_cnt_i0 (.D(n10374), .CK(clk_N_168), .CD(n18799), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[3] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_3), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_3), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[3] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15331), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15330), .COUT(n15331), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15329), .COUT(n15330), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15328), .COUT(n15329), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15327), .COUT(n15328), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15326), .COUT(n15327), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15325), .COUT(n15326), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15324), .COUT(n15325), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15323), .COUT(n15324), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15322), .COUT(n15323), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15321), .COUT(n15322), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15320), .COUT(n15321), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15319), .COUT(n15320), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15318), .COUT(n15319), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_351), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_356), .CD(n18799), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=74, LSE_RLINE=80 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15317), .COUT(n15318), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10225)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_768), .B(n58), .C(n52), .D(n40_adj_769), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_768)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_769)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12288_2_lut (.A(delay_cnt[0]), .B(n10225), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12288_2_lut.init = 16'h2222;
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15316), .COUT(n15317), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15316), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 key_reg_I_0_2_lut_rep_617 (.A(key_reg), .B(key_c_3), .Z(n18799)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_617.init = 16'h6666;
    LUT4 i7472_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7472_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7473_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7473_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7475_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7475_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7476_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7476_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7478_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7478_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7479_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7479_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_3), .C(n10225), .D(delay_cnt[0]), 
         .Z(clk_N_168_enable_351)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i7480_2_lut_3_lut (.A(key_reg), .B(key_c_3), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7480_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i5530_2_lut_rep_454 (.A(delay_cnt[0]), .B(n10225), .Z(clk_N_168_enable_356)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5530_2_lut_rep_454.init = 16'heeee;
    LUT4 i5531_2_lut_3_lut (.A(delay_cnt[0]), .B(n10225), .C(n9[0]), .Z(n10374)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5531_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_554 (.A(\key_flag[3] ), .B(\key_value[3] ), .Z(n18736)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_554.init = 16'h2222;
    LUT4 i285_3_lut_4_lut (.A(\key_flag[3] ), .B(\key_value[3] ), .C(n6), 
         .D(n18814), .Z(n887)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i285_3_lut_4_lut.init = 16'h2220;
    LUT4 n446_bdd_3_lut_4_lut (.A(\key_flag[3] ), .B(\key_value[3] ), .C(\rom2[1] ), 
         .D(n18754), .Z(n18598)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam n446_bdd_3_lut_4_lut.init = 16'hf202;
    LUT4 i1_2_lut_rep_525_3_lut_4_lut (.A(\key_flag[3] ), .B(\key_value[3] ), 
         .C(\key_flag[2] ), .D(\key_value[2] ), .Z(n18707)) /* synthesis lut_function=(!(A (B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_525_3_lut_4_lut.init = 16'h22f2;
    LUT4 i97_3_lut_4_lut (.A(\key_flag[3] ), .B(\key_value[3] ), .C(n18747), 
         .D(n18758), .Z(n444)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i97_3_lut_4_lut.init = 16'h2220;
    LUT4 i1_2_lut_rep_514_3_lut_4_lut (.A(\key_flag[3] ), .B(\key_value[3] ), 
         .C(\key_value[4] ), .D(\key_flag[4] ), .Z(n18696)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (C+!(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam i1_2_lut_rep_514_3_lut_4_lut.init = 16'h2f22;
    
endmodule
//
// Verilog Description of module clk_pll
//

module clk_pll (sys_clk_c, clk, GND_net, clk_N_168) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input sys_clk_c;
    output clk;
    input GND_net;
    output clk_N_168;
    
    wire sys_clk_c /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(3[12:19])
    wire clk /* synthesis is_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(13[7:10])
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    
    EHXPLLJ PLLInst_0 (.CLKI(sys_clk_c), .CLKFB(clk), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(clk)) /* synthesis FREQUENCY_PIN_CLKOP="48.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="8", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=1, LSE_LCOL=9, LSE_RCOL=5, LSE_LLINE=31, LSE_RLINE=34 */ ;   // d:/fpga_project/lattice_diamond/piano/piano.v(31[9] 34[5])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 4;
    defparam PLLInst_0.CLKOP_DIV = 11;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 10;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    INV i12987 (.A(clk), .Z(clk_N_168));
    
endmodule
//
// Verilog Description of module key_U23
//

module key_U23 (clk_N_168, \key_flag[13] , key_c_13, \key_value[13] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input clk_N_168;
    output \key_flag[13] ;
    input key_c_13;
    output \key_value[13] ;
    input GND_net;
    
    wire clk_N_168 /* synthesis is_inv_clock=1 */ ;   // d:/fpga_project/lattice_diamond/piano/speaker.v(16[13:21])
    wire [31:0]delay_cnt;   // d:/fpga_project/lattice_diamond/piano/key.v(12[13:22])
    
    wire n18789, n10394, key_flag_N_639, key_reg, clk_N_168_enable_46;
    wire [31:0]n9;
    
    wire clk_N_168_enable_41;
    wire [31:0]delay_cnt_31__N_570;
    
    wire n15560, n15559, n15558, n15557, n15556, n15555, n15554, 
        n15553, n15552, n15551, n15550, n15549, n15548, n15547, 
        n15546, n15545, n10258, n55, n60, n49, n50, n48, n39_adj_766, 
        n58, n52, n40_adj_767, n54, n44;
    
    FD1S3IX delay_cnt_i0 (.D(n10394), .CK(clk_N_168), .CD(n18789), .Q(delay_cnt[0])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i0.GSR = "ENABLED";
    FD1S3AX key_flag_27 (.D(key_flag_N_639), .CK(clk_N_168), .Q(\key_flag[13] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_flag_27.GSR = "ENABLED";
    FD1S3AY key_reg_25 (.D(key_c_13), .CK(clk_N_168), .Q(key_reg)) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam key_reg_25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i31 (.D(n9[31]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[31])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i31.GSR = "ENABLED";
    FD1P3IX delay_cnt_i30 (.D(n9[30]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[30])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i30.GSR = "ENABLED";
    FD1P3IX delay_cnt_i29 (.D(n9[29]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[29])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i29.GSR = "ENABLED";
    FD1P3IX delay_cnt_i28 (.D(n9[28]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[28])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i27 (.D(n9[27]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[27])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i27.GSR = "ENABLED";
    FD1P3IX delay_cnt_i26 (.D(n9[26]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[26])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i26.GSR = "ENABLED";
    FD1P3IX delay_cnt_i25 (.D(n9[25]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[25])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i25.GSR = "ENABLED";
    FD1P3IX delay_cnt_i24 (.D(n9[24]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[24])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i24.GSR = "ENABLED";
    FD1P3IX delay_cnt_i23 (.D(n9[23]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[23])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i23.GSR = "ENABLED";
    FD1P3IX delay_cnt_i22 (.D(n9[22]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[22])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i22.GSR = "ENABLED";
    FD1P3AX delay_cnt_i17 (.D(delay_cnt_31__N_570[17]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[17])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i17.GSR = "ENABLED";
    FD1P3AX delay_cnt_i18 (.D(delay_cnt_31__N_570[18]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[18])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i18.GSR = "ENABLED";
    FD1P3AX delay_cnt_i19 (.D(delay_cnt_31__N_570[19]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[19])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i19.GSR = "ENABLED";
    FD1P3IX delay_cnt_i20 (.D(n9[20]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[20])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i20.GSR = "ENABLED";
    FD1P3IX delay_cnt_i21 (.D(n9[21]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[21])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i21.GSR = "ENABLED";
    FD1P3AX delay_cnt_i16 (.D(delay_cnt_31__N_570[16]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[16])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i16.GSR = "ENABLED";
    FD1P3IX delay_cnt_i15 (.D(n9[15]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[15])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i15.GSR = "ENABLED";
    FD1P3AX delay_cnt_i14 (.D(delay_cnt_31__N_570[14]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[14])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i14.GSR = "ENABLED";
    FD1P3IX delay_cnt_i13 (.D(n9[13]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[13])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i13.GSR = "ENABLED";
    FD1P3IX delay_cnt_i12 (.D(n9[12]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[12])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i12.GSR = "ENABLED";
    FD1P3IX delay_cnt_i11 (.D(n9[11]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[11])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i11.GSR = "ENABLED";
    FD1P3IX delay_cnt_i10 (.D(n9[10]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[10])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i10.GSR = "ENABLED";
    FD1P3AX delay_cnt_i9 (.D(delay_cnt_31__N_570[9]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[9])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i9.GSR = "ENABLED";
    FD1P3AY key_value_28 (.D(key_c_13), .SP(key_flag_N_639), .CK(clk_N_168), 
            .Q(\key_value[13] )) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(38[18] 47[14])
    defparam key_value_28.GSR = "ENABLED";
    FD1P3IX delay_cnt_i8 (.D(n9[8]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[8])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i8.GSR = "ENABLED";
    FD1P3IX delay_cnt_i7 (.D(n9[7]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[7])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i7.GSR = "ENABLED";
    FD1P3AX delay_cnt_i6 (.D(delay_cnt_31__N_570[6]), .SP(clk_N_168_enable_41), 
            .CK(clk_N_168), .Q(delay_cnt[6])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i6.GSR = "ENABLED";
    FD1P3IX delay_cnt_i5 (.D(n9[5]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[5])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i5.GSR = "ENABLED";
    FD1P3IX delay_cnt_i4 (.D(n9[4]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[4])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i4.GSR = "ENABLED";
    FD1P3IX delay_cnt_i3 (.D(n9[3]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[3])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i3.GSR = "ENABLED";
    FD1P3IX delay_cnt_i2 (.D(n9[2]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[2])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i2.GSR = "ENABLED";
    FD1P3IX delay_cnt_i1 (.D(n9[1]), .SP(clk_N_168_enable_46), .CD(n18789), 
            .CK(clk_N_168), .Q(delay_cnt[1])) /* synthesis LSE_LINE_FILE_ID=1, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=156, LSE_RLINE=162 */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(20[16] 30[15])
    defparam delay_cnt_i1.GSR = "ENABLED";
    CCU2D sub_10_add_2_33 (.A0(delay_cnt[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n15560), .S0(n9[31]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_33.INIT0 = 16'h5555;
    defparam sub_10_add_2_33.INIT1 = 16'h0000;
    defparam sub_10_add_2_33.INJECT1_0 = "NO";
    defparam sub_10_add_2_33.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_31 (.A0(delay_cnt[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15559), .COUT(n15560), .S0(n9[29]), .S1(n9[30]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_31.INIT0 = 16'h5555;
    defparam sub_10_add_2_31.INIT1 = 16'h5555;
    defparam sub_10_add_2_31.INJECT1_0 = "NO";
    defparam sub_10_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_29 (.A0(delay_cnt[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15558), .COUT(n15559), .S0(n9[27]), .S1(n9[28]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_29.INIT0 = 16'h5555;
    defparam sub_10_add_2_29.INIT1 = 16'h5555;
    defparam sub_10_add_2_29.INJECT1_0 = "NO";
    defparam sub_10_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_27 (.A0(delay_cnt[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15557), .COUT(n15558), .S0(n9[25]), .S1(n9[26]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_27.INIT0 = 16'h5555;
    defparam sub_10_add_2_27.INIT1 = 16'h5555;
    defparam sub_10_add_2_27.INJECT1_0 = "NO";
    defparam sub_10_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_25 (.A0(delay_cnt[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15556), .COUT(n15557), .S0(n9[23]), .S1(n9[24]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_25.INIT0 = 16'h5555;
    defparam sub_10_add_2_25.INIT1 = 16'h5555;
    defparam sub_10_add_2_25.INJECT1_0 = "NO";
    defparam sub_10_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_23 (.A0(delay_cnt[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15555), .COUT(n15556), .S0(n9[21]), .S1(n9[22]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_23.INIT0 = 16'h5555;
    defparam sub_10_add_2_23.INIT1 = 16'h5555;
    defparam sub_10_add_2_23.INJECT1_0 = "NO";
    defparam sub_10_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_21 (.A0(delay_cnt[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15554), .COUT(n15555), .S0(n9[19]), .S1(n9[20]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_21.INIT0 = 16'h5555;
    defparam sub_10_add_2_21.INIT1 = 16'h5555;
    defparam sub_10_add_2_21.INJECT1_0 = "NO";
    defparam sub_10_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_19 (.A0(delay_cnt[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15553), .COUT(n15554), .S0(n9[17]), .S1(n9[18]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_19.INIT0 = 16'h5555;
    defparam sub_10_add_2_19.INIT1 = 16'h5555;
    defparam sub_10_add_2_19.INJECT1_0 = "NO";
    defparam sub_10_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_17 (.A0(delay_cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15552), .COUT(n15553), .S0(n9[15]), .S1(n9[16]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h5555;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(delay_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15551), .COUT(n15552), .S0(n9[13]), .S1(n9[14]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_13 (.A0(delay_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15550), .COUT(n15551), .S0(n9[11]), .S1(n9[12]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(delay_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15549), .COUT(n15550), .S0(n9[9]), .S1(n9[10]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(delay_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15548), .COUT(n15549), .S0(n9[7]), .S1(n9[8]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(delay_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15547), .COUT(n15548), .S0(n9[5]), .S1(n9[6]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(delay_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15546), .COUT(n15547), .S0(n9[3]), .S1(n9[4]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(delay_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(delay_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n15545), .COUT(n15546), .S0(n9[1]), .S1(n9[2]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(delay_cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n15545), .S1(n9[0]));   // d:/fpga_project/lattice_diamond/piano/key.v(26[31:47])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i5550_2_lut_rep_443 (.A(delay_cnt[0]), .B(n10258), .Z(clk_N_168_enable_46)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5550_2_lut_rep_443.init = 16'heeee;
    LUT4 i5551_2_lut_3_lut (.A(delay_cnt[0]), .B(n10258), .C(n9[0]), .Z(n10394)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(28[19:42])
    defparam i5551_2_lut_3_lut.init = 16'he0e0;
    LUT4 key_reg_I_0_2_lut_rep_607 (.A(key_reg), .B(key_c_13), .Z(n18789)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam key_reg_I_0_2_lut_rep_607.init = 16'h6666;
    LUT4 i7342_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[14]), .Z(delay_cnt_31__N_570[14])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7342_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7341_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[16]), .Z(delay_cnt_31__N_570[16])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7341_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7338_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[19]), .Z(delay_cnt_31__N_570[19])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7338_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7339_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[18]), .Z(delay_cnt_31__N_570[18])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7339_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7340_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[17]), .Z(delay_cnt_31__N_570[17])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7340_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7343_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[9]), .Z(delay_cnt_31__N_570[9])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7343_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i7344_2_lut_3_lut (.A(key_reg), .B(key_c_13), .C(n9[6]), .Z(delay_cnt_31__N_570[6])) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i7344_2_lut_3_lut.init = 16'hf6f6;
    LUT4 i1_2_lut_3_lut_4_lut (.A(key_reg), .B(key_c_13), .C(n10258), 
         .D(delay_cnt[0]), .Z(clk_N_168_enable_41)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(24[24:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff6;
    LUT4 i30_4_lut (.A(n55), .B(n60), .C(n49), .D(n50), .Z(n10258)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i30_4_lut.init = 16'hfffe;
    LUT4 i24_4_lut (.A(delay_cnt[15]), .B(n48), .C(delay_cnt[31]), .D(delay_cnt[3]), 
         .Z(n55)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i24_4_lut.init = 16'hfffe;
    LUT4 i29_4_lut (.A(n39_adj_766), .B(n58), .C(n52), .D(n40_adj_767), 
         .Z(n60)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i29_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(delay_cnt[22]), .B(delay_cnt[28]), .C(delay_cnt[26]), 
         .D(delay_cnt[10]), .Z(n49)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i19_4_lut (.A(delay_cnt[17]), .B(delay_cnt[1]), .C(delay_cnt[18]), 
         .D(delay_cnt[2]), .Z(n50)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i17_4_lut (.A(delay_cnt[20]), .B(delay_cnt[16]), .C(delay_cnt[4]), 
         .D(delay_cnt[13]), .Z(n48)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i8_2_lut (.A(delay_cnt[8]), .B(delay_cnt[29]), .Z(n39_adj_766)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i8_2_lut.init = 16'heeee;
    LUT4 i27_4_lut (.A(delay_cnt[9]), .B(n54), .C(n44), .D(delay_cnt[12]), 
         .Z(n58)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i27_4_lut.init = 16'hfffe;
    LUT4 i21_4_lut (.A(delay_cnt[19]), .B(delay_cnt[25]), .C(delay_cnt[21]), 
         .D(delay_cnt[6]), .Z(n52)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i21_4_lut.init = 16'hfffe;
    LUT4 i9_2_lut (.A(delay_cnt[7]), .B(delay_cnt[11]), .Z(n40_adj_767)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i9_2_lut.init = 16'heeee;
    LUT4 i23_4_lut (.A(delay_cnt[27]), .B(delay_cnt[14]), .C(delay_cnt[30]), 
         .D(delay_cnt[5]), .Z(n54)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i23_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut (.A(delay_cnt[24]), .B(delay_cnt[23]), .Z(n44)) /* synthesis lut_function=(A+(B)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i13_2_lut.init = 16'heeee;
    LUT4 i12320_2_lut (.A(delay_cnt[0]), .B(n10258), .Z(key_flag_N_639)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/fpga_project/lattice_diamond/piano/key.v(39[16:34])
    defparam i12320_2_lut.init = 16'h2222;
    
endmodule
